** Name: two_stage_single_output_op_amp_122_11

.MACRO two_stage_single_output_op_amp_122_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=2e-6 W=10e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=47e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=221e-6
mTelescopicFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=264e-6
mMainBias5 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=11e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mTelescopicFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=8e-6 W=23e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=23e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=23e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=453e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=221e-6
mSecondStage1StageBias13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=474e-6
mTelescopicFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=8e-6 W=23e-6
mMainBias15 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=260e-6
mTelescopicFirstStageStageBias17 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=264e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=24e-6
mTelescopicFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=24e-6
mTelescopicFirstStageLoad20 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=148e-6
mMainBias22 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=55e-6
mSecondStage1Transconductor23 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=598e-6
mTelescopicFirstStageLoad24 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=10e-6
mMainBias25 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=58e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_122_11

** Expected Performance Values: 
** Gain: 190 dB
** Power consumption: 4.16401 mW
** Area: 13899 (mu_m)^2
** Transit frequency: 2.57701 MHz
** Transit frequency with error factor: 2.57728 MHz
** Slew rate: 12.3916 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 4.21001 V
** VoutMin: 0.710001 V
** VcmMax: 5.03001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 9.00701e+06 muA
** NormalTransistorNmos: 2.59758e+08 muA
** NormalTransistorPmos: -4.67709e+07 muA
** NormalTransistorPmos: -4.49179e+07 muA
** NormalTransistorNmos: 5.47601e+06 muA
** NormalTransistorNmos: 5.47601e+06 muA
** NormalTransistorPmos: -5.47699e+06 muA
** NormalTransistorPmos: -5.47799e+06 muA
** NormalTransistorPmos: -5.47699e+06 muA
** NormalTransistorPmos: -5.47799e+06 muA
** NormalTransistorNmos: 5.58701e+07 muA
** DiodeTransistorNmos: 5.58701e+07 muA
** NormalTransistorNmos: 5.47601e+06 muA
** NormalTransistorNmos: 5.47601e+06 muA
** NormalTransistorNmos: 4.51398e+08 muA
** NormalTransistorNmos: 4.51397e+08 muA
** NormalTransistorPmos: -4.51397e+08 muA
** NormalTransistorPmos: -4.51398e+08 muA
** DiodeTransistorNmos: 4.67701e+07 muA
** NormalTransistorNmos: 4.67701e+07 muA
** DiodeTransistorNmos: 4.49171e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.00799e+06 muA
** DiodeTransistorPmos: -2.59757e+08 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 2.65001  V
** out: 2.5  V
** outFirstStage: 3.85001  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX3: 0.558001  V
** outVoltageBiasXXpXX0: 4.01001  V
** outVoltageBiasXXpXX1: 3.64501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.38401  V
** innerTransistorStack2Load2: 4.38401  V
** out1: 4.20901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.561001  V
** innerTransconductance: 4.41401  V
** inner: 0.555001  V


.END