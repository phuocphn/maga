** Name: two_stage_single_output_op_amp_8_10

.MACRO two_stage_single_output_op_amp_8_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=124e-6
mSecondStage1StageBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mSimpleFirstStageTransconductor4 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=92e-6
mSimpleFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=84e-6
mSecondStage1StageBias6 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSimpleFirstStageTransconductor7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=92e-6
mMainBias8 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=214e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=559e-6
mSecondStage1Transconductor10 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=124e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.5e-12
.EOM two_stage_single_output_op_amp_8_10

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 4.54301 mW
** Area: 5568 (mu_m)^2
** Transit frequency: 7.00201 MHz
** Transit frequency with error factor: 6.99306 MHz
** Slew rate: 7.17855 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** negPSRR: 167 dB
** posPSRR: 97 dB
** VoutMax: 4.52001 V
** VoutMin: 0.190001 V
** VcmMax: 4.60001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorNmos: 2.13221e+08 muA
** DiodeTransistorPmos: -4.14719e+07 muA
** NormalTransistorPmos: -4.14719e+07 muA
** NormalTransistorNmos: 8.29431e+07 muA
** NormalTransistorNmos: 4.14711e+07 muA
** NormalTransistorNmos: 4.14711e+07 muA
** NormalTransistorNmos: 6.0244e+08 muA
** NormalTransistorPmos: -6.02439e+08 muA
** NormalTransistorPmos: -6.0244e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.1322e+08 muA


** Expected Voltages: 
** ibias: 0.593001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.19001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.19801  V
** sourceTransconductance: 1.93201  V
** innerTransconductance: 4.48601  V


.END