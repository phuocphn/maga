** Name: two_stage_single_output_op_amp_57_9

.MACRO two_stage_single_output_op_amp_57_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=34e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=8e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=477e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=12e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=23e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=8e-6 W=32e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=59e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=59e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=34e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=477e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=8e-6 W=32e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=107e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=301e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=301e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=54e-6
mMainBias18 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=152e-6
mMainBias19 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=219e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=23e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.1001e-12
.EOM two_stage_single_output_op_amp_57_9

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 13.2281 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 5.33601 MHz
** Transit frequency with error factor: 5.33107 MHz
** Slew rate: 4.71325 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 1.87001 V
** VcmMax: 3.10001 V
** VcmMin: -0.109999 V


** Expected Currents: 
** NormalTransistorPmos: -1.54108e+08 muA
** NormalTransistorPmos: -2.60289e+07 muA
** NormalTransistorNmos: 7.59401e+07 muA
** NormalTransistorNmos: 1.30185e+08 muA
** NormalTransistorNmos: 7.59381e+07 muA
** NormalTransistorNmos: 1.30181e+08 muA
** DiodeTransistorPmos: -7.59389e+07 muA
** NormalTransistorPmos: -7.59389e+07 muA
** NormalTransistorPmos: -1.08485e+08 muA
** NormalTransistorPmos: -1.08484e+08 muA
** NormalTransistorPmos: -5.42429e+07 muA
** NormalTransistorPmos: -5.42429e+07 muA
** NormalTransistorNmos: 2.18507e+09 muA
** DiodeTransistorNmos: 2.18507e+09 muA
** NormalTransistorPmos: -2.18506e+09 muA
** DiodeTransistorNmos: 1.54109e+08 muA
** NormalTransistorNmos: 1.54108e+08 muA
** DiodeTransistorNmos: 2.60281e+07 muA
** DiodeTransistorNmos: 2.60271e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.27401  V
** inputVoltageBiasXXnXX2: 1.69801  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 1.13701  V
** outSourceVoltageBiasXXnXX2: 0.860001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.29601  V
** out1: 3.68801  V
** sourceGCC1: 0.818001  V
** sourceGCC2: 0.818001  V
** sourceTransconductance: 3.26401  V
** inner: 1.13401  V


.END