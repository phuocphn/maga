** Name: two_stage_single_output_op_amp_25_4

.MACRO two_stage_single_output_op_amp_25_4 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=26e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=26e-6
mSecondStage1StageBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=78e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=22e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=26e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=123e-6
mSecondStage1Transconductor8 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=460e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=26e-6
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=49e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=31e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=397e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=556e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=49e-6
mMainBias16 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=594e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.30001e-12
.EOM two_stage_single_output_op_amp_25_4

** Expected Performance Values: 
** Gain: 141 dB
** Power consumption: 5.21301 mW
** Area: 5711 (mu_m)^2
** Transit frequency: 3.42801 MHz
** Transit frequency with error factor: 3.42466 MHz
** Slew rate: 3.87769 V/mu_s
** Phase margin: 60.1606°
** CMRR: 104 dB
** negPSRR: 103 dB
** posPSRR: 112 dB
** VoutMax: 4 V
** VoutMin: 0.670001 V
** VcmMax: 3.23001 V
** VcmMin: 0.620001 V


** Expected Currents: 
** NormalTransistorPmos: -5.91649e+08 muA
** DiodeTransistorNmos: 1.41941e+07 muA
** NormalTransistorNmos: 1.41931e+07 muA
** NormalTransistorNmos: 1.41941e+07 muA
** DiodeTransistorNmos: 1.41931e+07 muA
** NormalTransistorPmos: -2.83889e+07 muA
** NormalTransistorPmos: -2.83879e+07 muA
** NormalTransistorPmos: -1.41949e+07 muA
** NormalTransistorPmos: -1.41949e+07 muA
** NormalTransistorNmos: 4.0251e+08 muA
** NormalTransistorNmos: 4.02509e+08 muA
** NormalTransistorPmos: -4.02509e+08 muA
** NormalTransistorPmos: -4.02508e+08 muA
** DiodeTransistorNmos: 5.9165e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.843001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.07101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.617001  V
** innerStageBias: 4.26501  V
** innerTransistorStack1Load1: 0.616001  V
** out1: 1.18201  V
** sourceTransconductance: 3.24401  V
** innerStageBias: 4.24001  V
** innerTransconductance: 0.438001  V


.END