** Name: two_stage_single_output_op_amp_46_3

.MACRO two_stage_single_output_op_amp_46_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=18e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=16e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=40e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=23e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=39e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=89e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=89e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=426e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=31e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=39e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=32e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=82e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=82e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=44e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=512e-6
mSecondStage1StageBias19 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=572e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=16e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.20001e-12
.EOM two_stage_single_output_op_amp_46_3

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 3.26901 mW
** Area: 7178 (mu_m)^2
** Transit frequency: 2.80301 MHz
** Transit frequency with error factor: 2.80294 MHz
** Slew rate: 5.35944 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 4.47001 V
** VoutMin: 0.510001 V
** VcmMax: 3.85001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.03068e+08 muA
** NormalTransistorNmos: 1.53561e+07 muA
** NormalTransistorNmos: 2.79681e+07 muA
** NormalTransistorNmos: 4.23781e+07 muA
** NormalTransistorNmos: 2.79681e+07 muA
** NormalTransistorNmos: 4.23781e+07 muA
** DiodeTransistorPmos: -2.79689e+07 muA
** DiodeTransistorPmos: -2.79699e+07 muA
** NormalTransistorPmos: -2.79689e+07 muA
** NormalTransistorPmos: -2.79699e+07 muA
** NormalTransistorPmos: -2.88229e+07 muA
** NormalTransistorPmos: -1.44109e+07 muA
** NormalTransistorPmos: -1.44109e+07 muA
** NormalTransistorNmos: 3.40549e+08 muA
** NormalTransistorPmos: -3.40548e+08 muA
** NormalTransistorPmos: -3.40549e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.03067e+08 muA
** DiodeTransistorPmos: -1.53569e+07 muA


** Expected Voltages: 
** ibias: 1.12201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.917001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX2: 4.16401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.18501  V
** innerTransistorStack2Load2: 4.18301  V
** out1: 3.30701  V
** sourceGCC1: 0.532001  V
** sourceGCC2: 0.532001  V
** sourceTransconductance: 3.37701  V
** innerStageBias: 4.50701  V


.END