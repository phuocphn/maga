** Name: two_stage_single_output_op_amp_30_11

.MACRO two_stage_single_output_op_amp_30_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=6e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=166e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=190e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=124e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=10e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=70e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=190e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=399e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=166e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mSecondStage1StageBias13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=415e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=70e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=344e-6
mSecondStage1Transconductor17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=343e-6
mSimpleFirstStageLoad18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=124e-6
mMainBias19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=49e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10e-12
.EOM two_stage_single_output_op_amp_30_11

** Expected Performance Values: 
** Gain: 145 dB
** Power consumption: 3.73601 mW
** Area: 14991 (mu_m)^2
** Transit frequency: 4.02201 MHz
** Transit frequency with error factor: 4.01711 MHz
** Slew rate: 3.79052 V/mu_s
** Phase margin: 60.1606°
** CMRR: 100 dB
** negPSRR: 178 dB
** posPSRR: 98 dB
** VoutMax: 4.59001 V
** VoutMin: 0.710001 V
** VcmMax: 4.63001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 6.67101e+06 muA
** NormalTransistorNmos: 3.95982e+08 muA
** NormalTransistorPmos: -3.29969e+07 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** DiodeTransistorNmos: 3.80921e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 2.63475e+08 muA
** NormalTransistorNmos: 2.63474e+08 muA
** NormalTransistorPmos: -2.63474e+08 muA
** NormalTransistorPmos: -2.63475e+08 muA
** DiodeTransistorNmos: 3.29961e+07 muA
** NormalTransistorNmos: 3.29961e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -6.67199e+06 muA
** DiodeTransistorPmos: -3.95981e+08 muA


** Expected Voltages: 
** ibias: 1.20501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.82201  V
** out: 2.5  V
** outFirstStage: 4.22801  V
** outInputVoltageBiasXXnXX1: 1.11801  V
** outSourceVoltageBiasXXnXX1: 0.559001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.22801  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.650001  V
** innerTransconductance: 4.45701  V
** inner: 0.559001  V


.END