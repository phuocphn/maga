** Name: two_stage_single_output_op_amp_76_7

.MACRO two_stage_single_output_op_amp_76_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=34e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=132e-6
mMainBias3 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=43e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=89e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=63e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=34e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=63e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=89e-6
mSecondStage1StageBias13 out inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=297e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=70e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=80e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=469e-6
mMainBias19 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=245e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=171e-6
mFoldedCascodeFirstStageLoad21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=80e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=59e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_76_7

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 13.2071 mW
** Area: 4766 (mu_m)^2
** Transit frequency: 7.87001 MHz
** Transit frequency with error factor: 7.87019 MHz
** Slew rate: 7.15991 V/mu_s
** Phase margin: 65.8902°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 0.260001 V
** VcmMax: 5.17001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorPmos: -5.98179e+07 muA
** NormalTransistorPmos: -4.69434e+08 muA
** NormalTransistorPmos: -2.48399e+08 muA
** NormalTransistorPmos: -3.24899e+07 muA
** NormalTransistorPmos: -5.37349e+07 muA
** NormalTransistorPmos: -3.24899e+07 muA
** NormalTransistorPmos: -5.37349e+07 muA
** DiodeTransistorNmos: 3.24891e+07 muA
** NormalTransistorNmos: 3.24891e+07 muA
** NormalTransistorNmos: 3.24891e+07 muA
** NormalTransistorNmos: 4.24871e+07 muA
** DiodeTransistorNmos: 4.24861e+07 muA
** NormalTransistorNmos: 2.12441e+07 muA
** NormalTransistorNmos: 2.12441e+07 muA
** NormalTransistorNmos: 1.73624e+09 muA
** NormalTransistorPmos: -1.73623e+09 muA
** DiodeTransistorNmos: 5.98171e+07 muA
** NormalTransistorNmos: 5.98161e+07 muA
** DiodeTransistorNmos: 4.69435e+08 muA
** DiodeTransistorNmos: 2.484e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.950001  V
** inputVoltageBiasXXnXX3: 0.667001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.20801  V
** outSourceVoltageBiasXXnXX1: 0.604001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.11201  V
** sourceGCC2: 4.11201  V
** sourceTransconductance: 1.90501  V
** inner: 0.603001  V


.END