** Name: two_stage_single_output_op_amp_122_9

.MACRO two_stage_single_output_op_amp_122_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=5e-6 W=22e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=22e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=326e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=62e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=9e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=72e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=72e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=72e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=22e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=22e-6
mSecondStage1StageBias13 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=5e-6 W=600e-6
mTelescopicFirstStageLoad14 outFirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=72e-6
mMainBias15 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=28e-6
mTelescopicFirstStageStageBias17 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=326e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=63e-6
mTelescopicFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=63e-6
mTelescopicFirstStageLoad20 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=166e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=540e-6
mTelescopicFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=166e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=8e-6
mMainBias24 outVoltageBiasXXnXX3 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=76e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.3001e-12
.EOM two_stage_single_output_op_amp_122_9

** Expected Performance Values: 
** Gain: 154 dB
** Power consumption: 2.18801 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 2.79201 MHz
** Transit frequency with error factor: 2.79182 MHz
** Slew rate: 7.14812 V/mu_s
** Phase margin: 60.7336°
** CMRR: 141 dB
** VoutMax: 4.83001 V
** VoutMin: 0.730001 V
** VcmMax: 4.91001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 9.47501e+06 muA
** NormalTransistorNmos: 1.28781e+07 muA
** NormalTransistorPmos: -8.42299e+06 muA
** NormalTransistorPmos: -7.84699e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorPmos: -2.28579e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorPmos: -2.28579e+07 muA
** NormalTransistorNmos: 1.24183e+08 muA
** DiodeTransistorNmos: 1.24183e+08 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.72615e+08 muA
** DiodeTransistorNmos: 2.72614e+08 muA
** NormalTransistorPmos: -2.72614e+08 muA
** DiodeTransistorNmos: 8.42201e+06 muA
** NormalTransistorNmos: 8.42101e+06 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 7.84691e+07 muA
** DiodeTransistorPmos: -9.47599e+06 muA
** DiodeTransistorPmos: -1.28789e+07 muA


** Expected Voltages: 
** ibias: 1.13701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.26801  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.569001  V
** outVoltageBiasXXnXX3: 2.65001  V
** outVoltageBiasXXpXX0: 3.79701  V
** outVoltageBiasXXpXX1: 3.70401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.42001  V
** innerTransistorStack2Load2: 4.42001  V
** out1: 4.08601  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.554001  V
** inner: 0.568001  V


.END