** Name: two_stage_single_output_op_amp_43_12

.MACRO two_stage_single_output_op_amp_43_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=10e-6 W=20e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=20e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=122e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=71e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=59e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=22e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=10e-6 W=13e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=90e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=90e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=122e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=10e-6 W=13e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=89e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=40e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=40e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=5e-6 W=370e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mMainBias19 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=346e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=393e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mMainBias22 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=590e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_43_12

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 5.11301 mW
** Area: 14642 (mu_m)^2
** Transit frequency: 5.31001 MHz
** Transit frequency with error factor: 5.30302 MHz
** Slew rate: 9.84316 V/mu_s
** Phase margin: 62.4525°
** CMRR: 93 dB
** VoutMax: 4.25 V
** VoutMin: 1.60001 V
** VcmMax: 3.80001 V
** VcmMin: -0.25 V


** Expected Currents: 
** NormalTransistorNmos: 7.44571e+07 muA
** NormalTransistorPmos: -9.92379e+07 muA
** NormalTransistorPmos: -5.90479e+07 muA
** NormalTransistorNmos: 4.44351e+07 muA
** NormalTransistorNmos: 7.61761e+07 muA
** NormalTransistorNmos: 4.44331e+07 muA
** NormalTransistorNmos: 7.61721e+07 muA
** DiodeTransistorPmos: -4.44339e+07 muA
** NormalTransistorPmos: -4.44339e+07 muA
** NormalTransistorPmos: -6.34789e+07 muA
** NormalTransistorPmos: -3.17399e+07 muA
** NormalTransistorPmos: -3.17399e+07 muA
** NormalTransistorNmos: 6.1745e+08 muA
** DiodeTransistorNmos: 6.17449e+08 muA
** NormalTransistorPmos: -6.17449e+08 muA
** NormalTransistorPmos: -6.1745e+08 muA
** DiodeTransistorNmos: 9.92371e+07 muA
** NormalTransistorNmos: 9.92381e+07 muA
** DiodeTransistorNmos: 5.90471e+07 muA
** DiodeTransistorNmos: 5.90461e+07 muA
** DiodeTransistorPmos: -7.44579e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.71301  V
** out: 2.5  V
** outFirstStage: 4.19701  V
** outInputVoltageBiasXXnXX1: 2.00201  V
** outSourceVoltageBiasXXnXX1: 1.00101  V
** outSourceVoltageBiasXXnXX2: 0.720001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.19801  V
** sourceGCC1: 0.670001  V
** sourceGCC2: 0.670001  V
** sourceTransconductance: 3.48401  V
** innerTransconductance: 4.76101  V
** inner: 1.00201  V


.END