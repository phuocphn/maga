** Name: two_stage_single_output_op_amp_133_5

.MACRO two_stage_single_output_op_amp_133_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mSimpleFirstStageLoad2 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=176e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=165e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=442e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=83e-6
mSimpleFirstStageLoad7 FirstStageYinnerOutputLoad1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=420e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=530e-6
mSimpleFirstStageLoad9 outFirstStage ibias sourceNmos sourceNmos nmos4 L=3e-6 W=420e-6
mMainBias10 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=270e-6
mMainBias11 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=128e-6
mSimpleFirstStageTransconductor12 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=351e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=474e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=165e-6
mSecondStage1StageBias16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=442e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=176e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=351e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.8001e-12
.EOM two_stage_single_output_op_amp_133_5

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 13.8241 mW
** Area: 14864 (mu_m)^2
** Transit frequency: 10.2151 MHz
** Transit frequency with error factor: 10.1726 MHz
** Slew rate: 24.7884 V/mu_s
** Phase margin: 60.1606°
** CMRR: 70 dB
** VoutMax: 3.19001 V
** VoutMin: 0.150001 V
** VcmMax: 3.08001 V
** VcmMin: -0.339999 V


** Expected Currents: 
** NormalTransistorNmos: 3.78909e+08 muA
** NormalTransistorNmos: 1.81585e+08 muA
** DiodeTransistorPmos: -7.96299e+07 muA
** DiodeTransistorPmos: -7.96309e+07 muA
** NormalTransistorPmos: -7.96299e+07 muA
** NormalTransistorPmos: -7.96309e+07 muA
** NormalTransistorNmos: 5.8875e+08 muA
** NormalTransistorNmos: 5.8875e+08 muA
** NormalTransistorPmos: -1.01824e+09 muA
** NormalTransistorPmos: -5.09119e+08 muA
** NormalTransistorPmos: -5.09119e+08 muA
** NormalTransistorNmos: 1.01684e+09 muA
** NormalTransistorPmos: -1.01683e+09 muA
** DiodeTransistorPmos: -1.01683e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.78908e+08 muA
** NormalTransistorPmos: -3.78909e+08 muA
** DiodeTransistorPmos: -1.81584e+08 muA


** Expected Voltages: 
** ibias: 0.629001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.62401  V
** outSourceVoltageBiasXXpXX1: 3.81201  V
** outVoltageBiasXXpXX2: 3.83301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.04301  V
** innerSourceLoad1: 3.76601  V
** innerTransistorStack2Load1: 3.76601  V
** sourceTransconductance: 3.81401  V
** inner: 3.80601  V


.END