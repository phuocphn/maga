** Name: two_stage_single_output_op_amp_5_1

.MACRO two_stage_single_output_op_amp_5_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias2 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=33e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=51e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=51e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=51e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=190e-6
mSimpleFirstStageLoad7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=51e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=134e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=160e-6
mMainBias10 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=31e-6
mSecondStage1StageBias11 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=134e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_5_1

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 1.31601 mW
** Area: 3936 (mu_m)^2
** Transit frequency: 4.23301 MHz
** Transit frequency with error factor: 4.2293 MHz
** Slew rate: 5.40404 V/mu_s
** Phase margin: 60.1606°
** CMRR: 104 dB
** negPSRR: 105 dB
** posPSRR: 226 dB
** VoutMax: 4.82001 V
** VoutMin: 0.150001 V
** VcmMax: 4.05001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -9.57499e+06 muA
** NormalTransistorNmos: 2.47121e+07 muA
** NormalTransistorNmos: 2.47111e+07 muA
** NormalTransistorNmos: 2.47101e+07 muA
** NormalTransistorNmos: 2.47111e+07 muA
** NormalTransistorPmos: -4.94219e+07 muA
** NormalTransistorPmos: -2.47109e+07 muA
** NormalTransistorPmos: -2.47109e+07 muA
** NormalTransistorNmos: 1.84113e+08 muA
** NormalTransistorPmos: -1.84112e+08 muA
** DiodeTransistorNmos: 9.57401e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.707001  V
** out: 2.5  V
** outFirstStage: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.556001  V
** innerTransistorStack1Load1: 0.151001  V
** innerTransistorStack2Load1: 0.151001  V
** sourceTransconductance: 3.26701  V


.END