** Name: two_stage_single_output_op_amp_36_12

.MACRO two_stage_single_output_op_amp_36_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=194e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=195e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=295e-6
mSimpleFirstStageLoad5 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=211e-6
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=136e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=5e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mSimpleFirstStageTransconductor9 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=41e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=195e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=194e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias13 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mSecondStage1StageBias14 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=295e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=41e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=81e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=136e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=481e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=264e-6
mSimpleFirstStageLoad20 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=5e-6 W=211e-6
mMainBias21 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=19e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.40001e-12
.EOM two_stage_single_output_op_amp_36_12

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 4.19301 mW
** Area: 14998 (mu_m)^2
** Transit frequency: 6.39301 MHz
** Transit frequency with error factor: 6.38905 MHz
** Slew rate: 6.02515 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** negPSRR: 108 dB
** posPSRR: 101 dB
** VoutMax: 4.28001 V
** VoutMin: 0.930001 V
** VcmMax: 3.92001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00071e+07 muA
** NormalTransistorNmos: 1.62124e+08 muA
** NormalTransistorPmos: -3.85629e+07 muA
** DiodeTransistorPmos: -1.95239e+07 muA
** DiodeTransistorPmos: -1.95249e+07 muA
** NormalTransistorPmos: -1.95239e+07 muA
** NormalTransistorPmos: -1.95249e+07 muA
** NormalTransistorNmos: 3.90451e+07 muA
** DiodeTransistorNmos: 3.90441e+07 muA
** NormalTransistorNmos: 1.95231e+07 muA
** NormalTransistorNmos: 1.95231e+07 muA
** NormalTransistorNmos: 5.7876e+08 muA
** DiodeTransistorNmos: 5.78761e+08 muA
** NormalTransistorPmos: -5.78759e+08 muA
** NormalTransistorPmos: -5.7876e+08 muA
** DiodeTransistorNmos: 3.85621e+07 muA
** NormalTransistorNmos: 3.85621e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.00079e+07 muA
** DiodeTransistorPmos: -1.62123e+08 muA


** Expected Voltages: 
** ibias: 1.33801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.06801  V
** outInputVoltageBiasXXnXX1: 1.11801  V
** outSourceVoltageBiasXXnXX1: 0.559001  V
** outSourceVoltageBiasXXnXX2: 0.670001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.51001  V
** innerSourceLoad1: 4.23501  V
** innerTransistorStack2Load1: 4.23501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.59901  V
** inner: 0.559001  V
** inner: 0.666001  V


.END