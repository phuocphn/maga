** Name: two_stage_single_output_op_amp_120_9

.MACRO two_stage_single_output_op_amp_120_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=43e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=102e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=285e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=12e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=5e-6 W=106e-6
mTelescopicFirstStageLoad7 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=198e-6
mMainBias8 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=402e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=38e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=86e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=86e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=43e-6
mMainBias13 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mSecondStage1StageBias15 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=285e-6
mTelescopicFirstStageLoad16 outFirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=38e-6
mTelescopicFirstStageStageBias17 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=102e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=5e-6 W=106e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=586e-6
mTelescopicFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=198e-6
mMainBias21 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=175e-6
mMainBias22 outVoltageBiasXXnXX3 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=158e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.5e-12
.EOM two_stage_single_output_op_amp_120_9

** Expected Performance Values: 
** Gain: 145 dB
** Power consumption: 3.56801 mW
** Area: 13472 (mu_m)^2
** Transit frequency: 3.07201 MHz
** Transit frequency with error factor: 3.07161 MHz
** Slew rate: 4.69467 V/mu_s
** Phase margin: 60.1606°
** CMRR: 152 dB
** VoutMax: 4.54001 V
** VoutMin: 0.840001 V
** VcmMax: 3.75 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 5.72261e+07 muA
** NormalTransistorPmos: -2.49629e+07 muA
** NormalTransistorPmos: -2.26309e+07 muA
** NormalTransistorNmos: 1.81991e+07 muA
** NormalTransistorNmos: 1.81991e+07 muA
** DiodeTransistorPmos: -1.81999e+07 muA
** DiodeTransistorPmos: -1.82009e+07 muA
** NormalTransistorPmos: -1.81999e+07 muA
** NormalTransistorPmos: -1.82009e+07 muA
** NormalTransistorNmos: 5.90291e+07 muA
** DiodeTransistorNmos: 5.90281e+07 muA
** NormalTransistorNmos: 1.82001e+07 muA
** NormalTransistorNmos: 1.82001e+07 muA
** NormalTransistorNmos: 5.62393e+08 muA
** DiodeTransistorNmos: 5.62394e+08 muA
** NormalTransistorPmos: -5.62392e+08 muA
** DiodeTransistorNmos: 2.49621e+07 muA
** NormalTransistorNmos: 2.49611e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 2.26301e+07 muA
** DiodeTransistorPmos: -5.72269e+07 muA


** Expected Voltages: 
** ibias: 1.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.25701  V
** out: 2.5  V
** outFirstStage: 3.97101  V
** outInputVoltageBiasXXnXX1: 1.24601  V
** outSourceVoltageBiasXXnXX1: 0.623001  V
** outSourceVoltageBiasXXnXX2: 0.622001  V
** outVoltageBiasXXnXX3: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.21601  V
** innerTransistorStack2Load2: 4.21501  V
** out1: 3.49101  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.621001  V
** inner: 0.619001  V


.END