** Name: two_stage_single_output_op_amp_59_8

.MACRO two_stage_single_output_op_amp_59_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=144e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=58e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=266e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 outInputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=134e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=25e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=25e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=275e-6
mSecondStage1StageBias10 out outInputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=342e-6
mFoldedCascodeFirstStageLoad11 outFirstStage outInputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=134e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=129e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=266e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=422e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=422e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=71e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=430e-6
mFoldedCascodeFirstStageLoad18 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=3e-6 W=317e-6
mMainBias19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=449e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.5e-12
.EOM two_stage_single_output_op_amp_59_8

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 14.9991 mW
** Area: 14826 (mu_m)^2
** Transit frequency: 5.48901 MHz
** Transit frequency with error factor: 5.48925 MHz
** Slew rate: 7.86733 V/mu_s
** Phase margin: 60.1606°
** CMRR: 136 dB
** VoutMax: 4.25 V
** VoutMin: 1.69001 V
** VcmMax: 3.09001 V
** VcmMin: 0.110001 V


** Expected Currents: 
** NormalTransistorPmos: -4.4691e+08 muA
** NormalTransistorNmos: 1.30794e+08 muA
** NormalTransistorNmos: 1.96189e+08 muA
** NormalTransistorNmos: 1.30795e+08 muA
** NormalTransistorNmos: 1.9619e+08 muA
** NormalTransistorPmos: -1.30793e+08 muA
** NormalTransistorPmos: -1.30794e+08 muA
** DiodeTransistorPmos: -1.30793e+08 muA
** NormalTransistorPmos: -1.3079e+08 muA
** NormalTransistorPmos: -1.30789e+08 muA
** NormalTransistorPmos: -6.53959e+07 muA
** NormalTransistorPmos: -6.53959e+07 muA
** NormalTransistorNmos: 2.14062e+09 muA
** NormalTransistorNmos: 2.14061e+09 muA
** NormalTransistorPmos: -2.14061e+09 muA
** DiodeTransistorNmos: 4.46913e+08 muA
** DiodeTransistorNmos: 4.46914e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.91501  V
** outSourceVoltageBiasXXnXX1: 1.08301  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.14801  V
** innerStageBias: 4.29301  V
** out1: 3.32201  V
** sourceGCC1: 1.26901  V
** sourceGCC2: 1.26901  V
** sourceTransconductance: 3.29101  V
** innerStageBias: 0.899001  V


.END