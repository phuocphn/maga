** Name: two_stage_single_output_op_amp_78_10

.MACRO two_stage_single_output_op_amp_78_10 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=10e-6 W=96e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=10e-6 W=96e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=20e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=30e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=572e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=10e-6 W=96e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=30e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=20e-6
mSecondStage1StageBias13 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=585e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=96e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=130e-6
mMainBias16 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=39e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerOutputLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=29e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=340e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=340e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=588e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=226e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=29e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=147e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_78_10

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 5.05501 mW
** Area: 14799 (mu_m)^2
** Transit frequency: 4.46401 MHz
** Transit frequency with error factor: 4.46401 MHz
** Slew rate: 4.20722 V/mu_s
** Phase margin: 76.2034°
** CMRR: 147 dB
** VoutMax: 4.32001 V
** VoutMin: 0.210001 V
** VcmMax: 5.25 V
** VcmMin: 1.42001 V


** Expected Currents: 
** NormalTransistorNmos: 1.62454e+08 muA
** NormalTransistorNmos: 4.80501e+07 muA
** NormalTransistorPmos: -1.25849e+07 muA
** NormalTransistorPmos: -1.90489e+07 muA
** NormalTransistorPmos: -2.85719e+07 muA
** NormalTransistorPmos: -1.90529e+07 muA
** NormalTransistorPmos: -2.85779e+07 muA
** DiodeTransistorNmos: 1.90501e+07 muA
** DiodeTransistorNmos: 1.90511e+07 muA
** NormalTransistorNmos: 1.90521e+07 muA
** NormalTransistorNmos: 1.90511e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** DiodeTransistorNmos: 1.90461e+07 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 7.20742e+08 muA
** NormalTransistorPmos: -7.20741e+08 muA
** NormalTransistorPmos: -7.20742e+08 muA
** DiodeTransistorNmos: 1.25841e+07 muA
** NormalTransistorNmos: 1.25831e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.62453e+08 muA
** DiodeTransistorPmos: -4.80509e+07 muA


** Expected Voltages: 
** ibias: 0.615001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.17301  V
** outInputVoltageBiasXXnXX1: 1.26601  V
** outSourceVoltageBiasXXnXX1: 0.633001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.28201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.11601  V
** innerTransistorStack1Load2: 0.558001  V
** innerTransistorStack2Load2: 0.558001  V
** sourceGCC1: 4.44101  V
** sourceGCC2: 4.44101  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.67101  V
** inner: 0.632001  V


.END