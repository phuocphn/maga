** Name: one_stage_single_output_op_amp47

.MACRO one_stage_single_output_op_amp47 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=5e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=52e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=431e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=431e-6
mMainBias8 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=28e-6
mMainBias9 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=14e-6
mFoldedCascodeFirstStageLoad10 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=52e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=373e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=96e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=96e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=92e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=92e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=82e-6
mFoldedCascodeFirstStageLoad17 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=373e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp47

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 2.20201 mW
** Area: 7106 (mu_m)^2
** Transit frequency: 5.32401 MHz
** Transit frequency with error factor: 5.3242 MHz
** Slew rate: 6.79626 V/mu_s
** Phase margin: 87.0896°
** CMRR: 134 dB
** VoutMax: 4.47001 V
** VoutMin: 0.910001 V
** VcmMax: 3.62001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 6.66701e+06 muA
** NormalTransistorNmos: 1.3654e+08 muA
** NormalTransistorNmos: 2.05225e+08 muA
** NormalTransistorNmos: 1.3654e+08 muA
** NormalTransistorNmos: 2.05225e+08 muA
** NormalTransistorPmos: -1.36539e+08 muA
** NormalTransistorPmos: -1.3654e+08 muA
** NormalTransistorPmos: -1.36539e+08 muA
** NormalTransistorPmos: -1.3654e+08 muA
** NormalTransistorPmos: -1.37372e+08 muA
** NormalTransistorPmos: -6.86859e+07 muA
** NormalTransistorPmos: -6.86859e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.33339e+07 muA
** DiodeTransistorPmos: -6.66799e+06 muA


** Expected Voltages: 
** ibias: 1.26601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** inputVoltageBiasXXpXX2: 3.82301  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.15301  V
** innerTransistorStack1Load2: 4.49701  V
** innerTransistorStack2Load2: 4.49701  V
** sourceGCC1: 0.507001  V
** sourceGCC2: 0.507001  V
** sourceTransconductance: 3.26801  V


.END