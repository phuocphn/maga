** Name: one_stage_single_output_op_amp89

.MACRO one_stage_single_output_op_amp89 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=12e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=45e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=9e-6 W=9e-6
mTelescopicFirstStageLoad5 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=109e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=87e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=87e-6
mTelescopicFirstStageLoad8 out inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=109e-6
mMainBias9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=18e-6
mTelescopicFirstStageLoad10 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=9e-6 W=160e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=66e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=66e-6
mMainBias13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=55e-6
mTelescopicFirstStageLoad14 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=9e-6 W=160e-6
mMainBias15 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=16e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=5e-6 W=394e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp89

** Expected Performance Values: 
** Gain: 95 dB
** Power consumption: 0.624001 mW
** Area: 7679 (mu_m)^2
** Transit frequency: 3.52101 MHz
** Transit frequency with error factor: 3.52064 MHz
** Slew rate: 4.42924 V/mu_s
** Phase margin: 60.1606°
** CMRR: 147 dB
** VoutMax: 4.20001 V
** VoutMin: 0.300001 V
** VcmMax: 4 V
** VcmMin: -0.0499999 V


** Expected Currents: 
** NormalTransistorNmos: 5.33201e+06 muA
** NormalTransistorPmos: -3.60999e+06 muA
** NormalTransistorPmos: -1.23129e+07 muA
** NormalTransistorPmos: -4.17819e+07 muA
** NormalTransistorPmos: -4.17839e+07 muA
** NormalTransistorNmos: 4.17811e+07 muA
** NormalTransistorNmos: 4.17821e+07 muA
** NormalTransistorNmos: 4.17831e+07 muA
** NormalTransistorNmos: 4.17821e+07 muA
** NormalTransistorPmos: -8.88979e+07 muA
** NormalTransistorPmos: -4.17829e+07 muA
** NormalTransistorPmos: -4.17829e+07 muA
** DiodeTransistorNmos: 3.60901e+06 muA
** DiodeTransistorNmos: 1.23121e+07 muA
** DiodeTransistorPmos: -5.33299e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outVoltageBiasXXnXX0: 0.562001  V
** outVoltageBiasXXpXX1: 2.13901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.25201  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 3.06401  V
** sourceGCC2: 3.06401  V


.END