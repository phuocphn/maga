** Name: one_stage_single_output_op_amp53

.MACRO one_stage_single_output_op_amp53 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=13e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=8e-6 W=30e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=13e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=59e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=59e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=73e-6
mMainBias10 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=55e-6
mFoldedCascodeFirstStageLoad11 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=30e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=187e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=102e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=102e-6
mFoldedCascodeFirstStageLoad15 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=187e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp53

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 1.51701 mW
** Area: 2311 (mu_m)^2
** Transit frequency: 2.90201 MHz
** Transit frequency with error factor: 2.90153 MHz
** Slew rate: 3.78724 V/mu_s
** Phase margin: 88.8085°
** CMRR: 133 dB
** VoutMax: 4.03001 V
** VoutMin: 1.64001 V
** VcmMax: 5.15001 V
** VcmMin: 0.790001 V


** Expected Currents: 
** NormalTransistorNmos: 6.12351e+07 muA
** NormalTransistorPmos: -7.59469e+07 muA
** NormalTransistorPmos: -1.16089e+08 muA
** NormalTransistorPmos: -7.59469e+07 muA
** NormalTransistorPmos: -1.16089e+08 muA
** DiodeTransistorNmos: 7.59461e+07 muA
** DiodeTransistorNmos: 7.59451e+07 muA
** NormalTransistorNmos: 7.59461e+07 muA
** NormalTransistorNmos: 7.59451e+07 muA
** NormalTransistorNmos: 8.02841e+07 muA
** NormalTransistorNmos: 4.01421e+07 muA
** NormalTransistorNmos: 4.01421e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.12359e+07 muA
** DiodeTransistorPmos: -6.12349e+07 muA


** Expected Voltages: 
** ibias: 0.567001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.18301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 1.14501  V
** innerTransistorStack2Load2: 1.14101  V
** out1: 2.03701  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.875  V


.END