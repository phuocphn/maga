** Name: two_stage_single_output_op_amp_115_12

.MACRO two_stage_single_output_op_amp_115_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=6e-6 W=14e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=22e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=572e-6
mMainBias4 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=34e-6
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=127e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=24e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mTelescopicFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=580e-6
mTelescopicFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=30e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=15e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=15e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=22e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=22e-6
mSecondStage1StageBias15 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=572e-6
mTelescopicFirstStageLoad16 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=30e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=113e-6
mTelescopicFirstStageStageBias18 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=147e-6
mTelescopicFirstStageLoad19 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=127e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=306e-6
mMainBias21 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=139e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=560e-6
mTelescopicFirstStageLoad23 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=11e-6
mMainBias24 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=429e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.7001e-12
.EOM two_stage_single_output_op_amp_115_12

** Expected Performance Values: 
** Gain: 177 dB
** Power consumption: 6.85401 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 3.62801 MHz
** Transit frequency with error factor: 3.62797 MHz
** Slew rate: 11.0929 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 3.80001 V
** VoutMin: 0.700001 V
** VcmMax: 4.15001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorNmos: 7.14801e+06 muA
** NormalTransistorNmos: 3.67171e+07 muA
** NormalTransistorPmos: -4.20279e+07 muA
** NormalTransistorPmos: -1.28233e+08 muA
** NormalTransistorNmos: 2.85711e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorPmos: -2.85719e+07 muA
** NormalTransistorPmos: -2.85709e+07 muA
** DiodeTransistorPmos: -2.85719e+07 muA
** NormalTransistorNmos: 1.85373e+08 muA
** NormalTransistorNmos: 1.85372e+08 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 1.08945e+09 muA
** DiodeTransistorNmos: 1.08945e+09 muA
** NormalTransistorPmos: -1.08944e+09 muA
** NormalTransistorPmos: -1.08944e+09 muA
** DiodeTransistorNmos: 4.20271e+07 muA
** NormalTransistorNmos: 4.20261e+07 muA
** DiodeTransistorNmos: 1.28234e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.14899e+06 muA
** DiodeTransistorPmos: -3.67179e+07 muA


** Expected Voltages: 
** ibias: 1.18501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11001  V
** inputVoltageBiasXXpXX0: 4.04701  V
** out: 2.5  V
** outFirstStage: 3.80201  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX3: 0.556001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX1: 3.18901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.27701  V
** innerStageBias: 0.480001  V
** out1: 3.33001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.32201  V
** inner: 0.555001  V


.END