** Name: two_stage_single_output_op_amp_46_6

.MACRO two_stage_single_output_op_amp_46_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=347e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=317e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=11e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=184e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=458e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=441e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=441e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=591e-6
mSecondStage1Transconductor12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=593e-6
mFoldedCascodeFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=458e-6
mMainBias14 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=35e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=347e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=51e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=51e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=595e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=45e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=184e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=317e-6
mMainBias23 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=56e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.7001e-12
.EOM two_stage_single_output_op_amp_46_6

** Expected Performance Values: 
** Gain: 169 dB
** Power consumption: 14.9771 mW
** Area: 7792 (mu_m)^2
** Transit frequency: 8.82401 MHz
** Transit frequency with error factor: 8.82416 MHz
** Slew rate: 28.3135 V/mu_s
** Phase margin: 67.6091°
** CMRR: 128 dB
** VoutMax: 3.26001 V
** VoutMin: 0.360001 V
** VcmMax: 3.53001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 6.72881e+07 muA
** NormalTransistorPmos: -5.69159e+07 muA
** NormalTransistorPmos: -4.57129e+07 muA
** NormalTransistorNmos: 5.36813e+08 muA
** NormalTransistorNmos: 8.39941e+08 muA
** NormalTransistorNmos: 5.36813e+08 muA
** NormalTransistorNmos: 8.39941e+08 muA
** DiodeTransistorPmos: -5.36812e+08 muA
** DiodeTransistorPmos: -5.36813e+08 muA
** NormalTransistorPmos: -5.36812e+08 muA
** NormalTransistorPmos: -5.36813e+08 muA
** NormalTransistorPmos: -6.06253e+08 muA
** NormalTransistorPmos: -3.03126e+08 muA
** NormalTransistorPmos: -3.03126e+08 muA
** NormalTransistorNmos: 1.12564e+09 muA
** NormalTransistorNmos: 1.12564e+09 muA
** NormalTransistorPmos: -1.12563e+09 muA
** DiodeTransistorPmos: -1.12563e+09 muA
** DiodeTransistorNmos: 5.69151e+07 muA
** DiodeTransistorNmos: 4.57121e+07 muA
** DiodeTransistorPmos: -6.72889e+07 muA
** NormalTransistorPmos: -6.72899e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.10001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.69601  V
** outSourceVoltageBiasXXpXX1: 3.84801  V
** outVoltageBiasXXnXX1: 0.921001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.14101  V
** innerTransistorStack2Load2: 4.13901  V
** out1: 3.26801  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.63801  V
** innerTransconductance: 0.304001  V
** inner: 3.84301  V


.END