** Name: two_stage_single_output_op_amp_138_3

.MACRO two_stage_single_output_op_amp_138_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=35e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=6e-6 W=10e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=6e-6 W=10e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mSimpleFirstStageLoad7 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=7e-6 W=139e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=149e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=149e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=129e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=162e-6
mSimpleFirstStageLoad12 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=139e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=103e-6
mSimpleFirstStageTransconductor14 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=77e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=6e-6 W=10e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=582e-6
mSecondStage1StageBias18 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=411e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=6e-6 W=10e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=77e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.80001e-12
.EOM two_stage_single_output_op_amp_138_3

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 4.16501 mW
** Area: 8816 (mu_m)^2
** Transit frequency: 3.65101 MHz
** Transit frequency with error factor: 3.64915 MHz
** Slew rate: 6.02876 V/mu_s
** Phase margin: 60.1606°
** CMRR: 85 dB
** VoutMax: 4.32001 V
** VoutMin: 0.320001 V
** VcmMax: 3.92001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 3.55351e+07 muA
** NormalTransistorNmos: 2.81681e+07 muA
** DiodeTransistorPmos: -1.69219e+07 muA
** NormalTransistorPmos: -1.69219e+07 muA
** NormalTransistorPmos: -1.69219e+07 muA
** DiodeTransistorPmos: -1.69219e+07 muA
** NormalTransistorNmos: 4.06761e+07 muA
** NormalTransistorNmos: 4.06771e+07 muA
** NormalTransistorNmos: 4.06761e+07 muA
** NormalTransistorNmos: 4.06771e+07 muA
** NormalTransistorPmos: -4.75109e+07 muA
** NormalTransistorPmos: -2.37549e+07 muA
** NormalTransistorPmos: -2.37549e+07 muA
** NormalTransistorNmos: 6.779e+08 muA
** NormalTransistorPmos: -6.77899e+08 muA
** NormalTransistorPmos: -6.779e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.55359e+07 muA
** DiodeTransistorPmos: -2.81689e+07 muA


** Expected Voltages: 
** ibias: 1.11401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.721001  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outVoltageBiasXXpXX2: 4.18101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.553001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.553001  V
** sourceTransconductance: 3.32601  V
** innerStageBias: 4.67801  V


.END