** Name: two_stage_single_output_op_amp_195_10

.MACRO two_stage_single_output_op_amp_195_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=32e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=16e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mMainBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=599e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=77e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=32e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=21e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=32e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=9e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=9e-6 W=65e-6
mMainBias11 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=202e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=346e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=16e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=9e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=140e-6
mSimpleFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=69e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=459e-6
mMainBias18 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=440e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=407e-6
mSimpleFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=69e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_195_10

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 8.44501 mW
** Area: 12513 (mu_m)^2
** Transit frequency: 3.16901 MHz
** Transit frequency with error factor: 3.14431 MHz
** Slew rate: 3.53049 V/mu_s
** Phase margin: 68.182°
** CMRR: 92 dB
** VoutMax: 4.49001 V
** VoutMin: 0.160001 V
** VcmMax: 4.83001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 1.08303e+08 muA
** NormalTransistorNmos: 1.54244e+08 muA
** NormalTransistorPmos: -8.81397e+08 muA
** DiodeTransistorNmos: 1.27942e+08 muA
** DiodeTransistorNmos: 1.27943e+08 muA
** NormalTransistorNmos: 1.27942e+08 muA
** NormalTransistorNmos: 1.27943e+08 muA
** NormalTransistorPmos: -1.35927e+08 muA
** NormalTransistorPmos: -1.35927e+08 muA
** NormalTransistorNmos: 1.59721e+07 muA
** NormalTransistorNmos: 1.59731e+07 muA
** NormalTransistorNmos: 7.98601e+06 muA
** NormalTransistorNmos: 7.98601e+06 muA
** NormalTransistorNmos: 2.63167e+08 muA
** NormalTransistorPmos: -2.63166e+08 muA
** NormalTransistorPmos: -2.63167e+08 muA
** DiodeTransistorNmos: 8.81398e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.08302e+08 muA
** DiodeTransistorPmos: -1.54243e+08 muA


** Expected Voltages: 
** ibias: 0.570001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.799001  V
** inputVoltageBiasXXpXX2: 3.85901  V
** out: 2.5  V
** outFirstStage: 4.25601  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.940001  V
** innerStageBias: 0.232001  V
** innerTransistorStack2Load1: 0.940001  V
** out1: 2.09501  V
** sourceTransconductance: 1.91701  V
** innerTransconductance: 4.57801  V


.END