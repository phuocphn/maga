** Name: two_stage_single_output_op_amp_45_5

.MACRO two_stage_single_output_op_amp_45_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=7e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=5e-6
mMainBias5 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=6e-6 W=9e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=5e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=228e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=50e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=210e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=210e-6
mMainBias11 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias12 inputVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
mSecondStage1Transconductor13 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=190e-6
mFoldedCascodeFirstStageLoad14 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=50e-6
mMainBias15 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=30e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=65e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=65e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=6e-6 W=78e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=228e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=578e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_45_5

** Expected Performance Values: 
** Gain: 117 dB
** Power consumption: 6.04301 mW
** Area: 8446 (mu_m)^2
** Transit frequency: 5.62001 MHz
** Transit frequency with error factor: 5.62024 MHz
** Slew rate: 19.8236 V/mu_s
** Phase margin: 64.7443°
** CMRR: 126 dB
** VoutMax: 3.11001 V
** VoutMin: 0.580001 V
** VcmMax: 3.25 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.96201e+07 muA
** NormalTransistorNmos: 1.00071e+07 muA
** NormalTransistorNmos: 1.06751e+07 muA
** NormalTransistorNmos: 9.15451e+07 muA
** NormalTransistorNmos: 1.37338e+08 muA
** NormalTransistorNmos: 9.15451e+07 muA
** NormalTransistorNmos: 1.37338e+08 muA
** DiodeTransistorPmos: -9.15459e+07 muA
** NormalTransistorPmos: -9.15459e+07 muA
** NormalTransistorPmos: -9.15459e+07 muA
** NormalTransistorPmos: -9.15869e+07 muA
** NormalTransistorPmos: -4.57929e+07 muA
** NormalTransistorPmos: -4.57929e+07 muA
** NormalTransistorNmos: 8.83609e+08 muA
** NormalTransistorPmos: -8.83608e+08 muA
** DiodeTransistorPmos: -8.83609e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.96209e+07 muA
** NormalTransistorPmos: -1.96219e+07 muA
** DiodeTransistorPmos: -1.00079e+07 muA
** DiodeTransistorPmos: -1.06759e+07 muA


** Expected Voltages: 
** ibias: 1.18701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.68601  V
** inputVoltageBiasXXpXX3: 3.80501  V
** out: 2.5  V
** outFirstStage: 0.982001  V
** outInputVoltageBiasXXpXX1: 2.55001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 3.77501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.46001  V
** out1: 4.09601  V
** sourceGCC1: 0.526001  V
** sourceGCC2: 0.526001  V
** sourceTransconductance: 3.62301  V
** inner: 3.77401  V


.END