** Name: one_stage_single_output_op_amp52

.MACRO one_stage_single_output_op_amp52 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=84e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=35e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=23e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=84e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=22e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=22e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=286e-6
mFoldedCascodeFirstStageLoad10 out inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=131e-6
mFoldedCascodeFirstStageLoad11 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=212e-6
mFoldedCascodeFirstStageLoad12 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=184e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=184e-6
mMainBias14 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=38e-6
mMainBias15 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mFoldedCascodeFirstStageLoad16 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=212e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp52

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 2.23101 mW
** Area: 3829 (mu_m)^2
** Transit frequency: 5.39501 MHz
** Transit frequency with error factor: 5.39529 MHz
** Slew rate: 6.19449 V/mu_s
** Phase margin: 88.2356°
** CMRR: 143 dB
** VoutMax: 4.02001 V
** VoutMin: 0.470001 V
** VcmMax: 5.17001 V
** VcmMin: 0.75 V


** Expected Currents: 
** NormalTransistorPmos: -3.79269e+07 muA
** NormalTransistorPmos: -1.52079e+07 muA
** NormalTransistorPmos: -1.24368e+08 muA
** NormalTransistorPmos: -1.86551e+08 muA
** NormalTransistorPmos: -1.24369e+08 muA
** NormalTransistorPmos: -1.86552e+08 muA
** DiodeTransistorNmos: 1.24369e+08 muA
** NormalTransistorNmos: 1.2437e+08 muA
** NormalTransistorNmos: 1.24369e+08 muA
** NormalTransistorNmos: 1.24368e+08 muA
** NormalTransistorNmos: 6.21841e+07 muA
** NormalTransistorNmos: 6.21841e+07 muA
** DiodeTransistorNmos: 3.79261e+07 muA
** DiodeTransistorNmos: 1.52071e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.07101  V
** inputVoltageBiasXXnXX2: 0.565001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.387001  V
** out1: 0.592001  V
** sourceGCC1: 4.22401  V
** sourceGCC2: 4.22401  V
** sourceTransconductance: 1.91201  V


.END