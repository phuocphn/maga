** Name: two_stage_single_output_op_amp_1_3

.MACRO two_stage_single_output_op_amp_1_3 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=79e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=536e-6
mSimpleFirstStageLoad7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=79e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=22e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=66e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=141e-6
mMainBias11 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mSecondStage1StageBias12 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=119e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=22e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_1_3

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 1.33401 mW
** Area: 5785 (mu_m)^2
** Transit frequency: 2.90301 MHz
** Transit frequency with error factor: 2.88793 MHz
** Slew rate: 5.23556 V/mu_s
** Phase margin: 68.755°
** CMRR: 87 dB
** negPSRR: 89 dB
** posPSRR: 218 dB
** VoutMax: 4.53001 V
** VoutMin: 0.150001 V
** VcmMax: 3.48001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 4.04481e+07 muA
** NormalTransistorPmos: -1.65949e+07 muA
** DiodeTransistorNmos: 3.04251e+07 muA
** NormalTransistorNmos: 3.04251e+07 muA
** NormalTransistorPmos: -6.08479e+07 muA
** NormalTransistorPmos: -3.04239e+07 muA
** NormalTransistorPmos: -3.04239e+07 muA
** NormalTransistorNmos: 1.29008e+08 muA
** NormalTransistorPmos: -1.29007e+08 muA
** NormalTransistorPmos: -1.29008e+08 muA
** DiodeTransistorNmos: 1.65941e+07 muA
** DiodeTransistorPmos: -4.04489e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.686001  V
** inputVoltageBiasXXpXX1: 3.95801  V
** out: 2.5  V
** outFirstStage: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.556001  V
** sourceTransconductance: 3.79701  V
** innerStageBias: 4.76801  V


.END