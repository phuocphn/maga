** Name: two_stage_single_output_op_amp_187_8

.MACRO two_stage_single_output_op_amp_187_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=19e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=17e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=272e-6
mSimpleFirstStageStageBias5 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=84e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=21e-6
mSimpleFirstStageLoad7 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=19e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=35e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mSecondStage1StageBias10 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=243e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=7e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=21e-6
mMainBias13 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=388e-6
mSimpleFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=155e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=346e-6
mSimpleFirstStageLoad16 outFirstStage outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=155e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10e-12
.EOM two_stage_single_output_op_amp_187_8

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 3.45801 mW
** Area: 6972 (mu_m)^2
** Transit frequency: 4.22401 MHz
** Transit frequency with error factor: 4.20691 MHz
** Slew rate: 3.98052 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** VoutMax: 4.78001 V
** VoutMin: 0.790001 V
** VcmMax: 5.21001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 1.84782e+08 muA
** NormalTransistorNmos: 8.41651e+07 muA
** NormalTransistorNmos: 8.41641e+07 muA
** DiodeTransistorNmos: 8.41651e+07 muA
** NormalTransistorPmos: -1.04163e+08 muA
** NormalTransistorPmos: -1.04163e+08 muA
** NormalTransistorNmos: 3.99971e+07 muA
** NormalTransistorNmos: 3.99981e+07 muA
** NormalTransistorNmos: 1.99991e+07 muA
** NormalTransistorNmos: 1.99991e+07 muA
** NormalTransistorNmos: 2.88581e+08 muA
** NormalTransistorNmos: 2.8858e+08 muA
** NormalTransistorPmos: -2.8858e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.84781e+08 muA


** Expected Voltages: 
** ibias: 1.12601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.21901  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 4.24201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.488001  V
** innerTransistorStack2Load1: 1.13201  V
** out1: 2.28701  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.483001  V


.END