** Name: two_stage_single_output_op_amp_82_6

.MACRO two_stage_single_output_op_amp_82_6 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=59e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=59e-6
mMainBias3 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=40e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=79e-6
mSecondStage1StageBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mMainBias6 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=15e-6
mMainBias7 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=14e-6
mSecondStage1StageBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=346e-6
mMainBias9 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=288e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=59e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=29e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=79e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=128e-6
mMainBias15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=40e-6
mMainBias16 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=600e-6
mSecondStage1Transconductor17 out outVoltageBiasXXnXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=594e-6
mFoldedCascodeFirstStageLoad18 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=59e-6
mMainBias19 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=93e-6
mFoldedCascodeFirstStageLoad20 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=28e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=49e-6
mFoldedCascodeFirstStageLoad22 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=49e-6
mMainBias23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=14e-6
mSecondStage1StageBias24 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=346e-6
mFoldedCascodeFirstStageLoad25 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=28e-6
mMainBias26 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=412e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_82_6

** Expected Performance Values: 
** Gain: 172 dB
** Power consumption: 5.10401 mW
** Area: 14658 (mu_m)^2
** Transit frequency: 4.44401 MHz
** Transit frequency with error factor: 4.44398 MHz
** Slew rate: 3.54452 V/mu_s
** Phase margin: 64.7443°
** CMRR: 146 dB
** VoutMax: 3.58001 V
** VoutMin: 0.660001 V
** VcmMax: 5.23001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 2.30111e+07 muA
** NormalTransistorNmos: 1.51453e+08 muA
** NormalTransistorPmos: -2.19051e+08 muA
** NormalTransistorPmos: -1.60539e+07 muA
** NormalTransistorPmos: -2.58279e+07 muA
** NormalTransistorPmos: -1.60539e+07 muA
** NormalTransistorPmos: -2.58279e+07 muA
** DiodeTransistorNmos: 1.60531e+07 muA
** NormalTransistorNmos: 1.60541e+07 muA
** NormalTransistorNmos: 1.60531e+07 muA
** DiodeTransistorNmos: 1.60541e+07 muA
** NormalTransistorNmos: 1.95461e+07 muA
** DiodeTransistorNmos: 1.95471e+07 muA
** NormalTransistorNmos: 9.77301e+06 muA
** NormalTransistorNmos: 9.77301e+06 muA
** NormalTransistorNmos: 5.65675e+08 muA
** NormalTransistorNmos: 5.65674e+08 muA
** NormalTransistorPmos: -5.65674e+08 muA
** DiodeTransistorPmos: -5.65675e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 2.19052e+08 muA
** DiodeTransistorPmos: -2.30119e+07 muA
** NormalTransistorPmos: -2.30129e+07 muA
** DiodeTransistorPmos: -1.51452e+08 muA
** DiodeTransistorPmos: -1.51453e+08 muA


** Expected Voltages: 
** ibias: 1.13501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.95001  V
** out: 2.5  V
** outFirstStage: 0.915001  V
** outInputVoltageBiasXXpXX1: 3.01401  V
** outSourceVoltageBiasXXnXX1: 0.568001  V
** outSourceVoltageBiasXXpXX1: 4.00701  V
** outSourceVoltageBiasXXpXX2: 4.26401  V
** outVoltageBiasXXnXX2: 1.06501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.554001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.12001  V
** sourceGCC1: 3.69301  V
** sourceGCC2: 3.69301  V
** sourceTransconductance: 1.94001  V
** innerTransconductance: 0.510001  V
** inner: 0.567001  V
** inner: 4.00501  V


.END