** Name: two_stage_single_output_op_amp_76_2

.MACRO two_stage_single_output_op_amp_76_2 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=26e-6
mMainBias2 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=29e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=385e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=26e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=134e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=134e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=385e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=197e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=29e-6
mSecondStage1Transconductor13 out inputVoltageBiasXXnXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=286e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=99e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=503e-6
mMainBias16 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=220e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=209e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=78e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=78e-6
mMainBias20 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
mSecondStage1StageBias21 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=316e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=209e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.1001e-12
.EOM two_stage_single_output_op_amp_76_2

** Expected Performance Values: 
** Gain: 134 dB
** Power consumption: 7.44701 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 9.55301 MHz
** Transit frequency with error factor: 9.55294 MHz
** Slew rate: 12.2638 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 4.63001 V
** VoutMin: 0.470001 V
** VcmMax: 5.04001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 1.72607e+08 muA
** NormalTransistorNmos: 7.57771e+07 muA
** NormalTransistorPmos: -7.82229e+07 muA
** NormalTransistorPmos: -1.2484e+08 muA
** NormalTransistorPmos: -1.90667e+08 muA
** NormalTransistorPmos: -1.2484e+08 muA
** NormalTransistorPmos: -1.90667e+08 muA
** DiodeTransistorNmos: 1.24841e+08 muA
** NormalTransistorNmos: 1.24841e+08 muA
** NormalTransistorNmos: 1.24841e+08 muA
** NormalTransistorNmos: 1.31657e+08 muA
** DiodeTransistorNmos: 1.31658e+08 muA
** NormalTransistorNmos: 6.58281e+07 muA
** NormalTransistorNmos: 6.58281e+07 muA
** NormalTransistorNmos: 7.71412e+08 muA
** NormalTransistorNmos: 7.71411e+08 muA
** NormalTransistorPmos: -7.71411e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 7.82221e+07 muA
** DiodeTransistorPmos: -1.72606e+08 muA
** DiodeTransistorPmos: -7.57779e+07 muA


** Expected Voltages: 
** ibias: 1.14701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.01401  V
** out: 2.5  V
** outFirstStage: 0.619001  V
** outSourceVoltageBiasXXnXX1: 0.574001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.06801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.437001  V
** out1: 0.642001  V
** sourceGCC1: 4.43201  V
** sourceGCC2: 4.43201  V
** sourceTransconductance: 1.87901  V
** innerTransconductance: 0.356001  V
** inner: 0.573001  V


.END