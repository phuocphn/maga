** Name: one_stage_single_output_op_amp107

.MACRO one_stage_single_output_op_amp107 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=24e-6
mMainBias4 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=95e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=476e-6
mTelescopicFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=476e-6
mTelescopicFirstStageLoad9 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=95e-6
mMainBias10 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
mTelescopicFirstStageLoad11 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=226e-6
mTelescopicFirstStageStageBias12 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=252e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=8e-6 W=174e-6
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=8e-6 W=174e-6
mTelescopicFirstStageLoad15 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=226e-6
mMainBias16 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mMainBias17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mTelescopicFirstStageStageBias18 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=600e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp107

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 1.60901 mW
** Area: 14250 (mu_m)^2
** Transit frequency: 2.98401 MHz
** Transit frequency with error factor: 2.9837 MHz
** Slew rate: 12.6216 V/mu_s
** Phase margin: 88.8085°
** CMRR: 142 dB
** VoutMax: 3.41001 V
** VoutMin: 0.300001 V
** VcmMax: 3 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 7.11061e+07 muA
** NormalTransistorPmos: -2.12909e+07 muA
** NormalTransistorPmos: -2.69349e+07 muA
** NormalTransistorPmos: -9.12109e+07 muA
** NormalTransistorPmos: -9.12109e+07 muA
** NormalTransistorNmos: 9.12101e+07 muA
** NormalTransistorNmos: 9.12091e+07 muA
** NormalTransistorNmos: 9.12101e+07 muA
** NormalTransistorNmos: 9.12091e+07 muA
** NormalTransistorPmos: -2.53525e+08 muA
** NormalTransistorPmos: -2.53526e+08 muA
** NormalTransistorPmos: -9.12099e+07 muA
** NormalTransistorPmos: -9.12099e+07 muA
** DiodeTransistorNmos: 2.12901e+07 muA
** DiodeTransistorNmos: 2.69341e+07 muA
** DiodeTransistorPmos: -7.11069e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.48201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.655001  V
** outVoltageBiasXXnXX1: 0.705001  V
** outVoltageBiasXXpXX1: 2.34901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.54601  V
** innerSourceLoad2: 0.555001  V
** innerStageBias: 4.19901  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 3.06301  V
** sourceGCC2: 3.06301  V


.END