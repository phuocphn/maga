** Name: two_stage_single_output_op_amp_100_5

.MACRO two_stage_single_output_op_amp_100_5 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=39e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=285e-6
mMainBias3 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=1e-6 W=16e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=56e-6
mTelescopicFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=510e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mMainBias7 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=7e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=596e-6
mTelescopicFirstStageLoad9 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=39e-6
mMainBias10 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=46e-6
mMainBias11 outVoltageBiasXXpXX3 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=163e-6
mTelescopicFirstStageLoad12 FirstStageYout1 outVoltageBiasXXpXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=8e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=238e-6
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=238e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=56e-6
mMainBias16 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mMainBias17 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=274e-6
mSecondStage1StageBias18 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=600e-6
mTelescopicFirstStageLoad19 outFirstStage outVoltageBiasXXpXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=8e-6
mTelescopicFirstStageStageBias20 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=510e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.7001e-12
.EOM two_stage_single_output_op_amp_100_5

** Expected Performance Values: 
** Gain: 104 dB
** Power consumption: 4.24501 mW
** Area: 11285 (mu_m)^2
** Transit frequency: 4.29101 MHz
** Transit frequency with error factor: 4.28754 MHz
** Slew rate: 9.71454 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** VoutMax: 4.06001 V
** VoutMin: 0.150001 V
** VcmMax: 3 V
** VcmMin: 1.91001 V


** Expected Currents: 
** NormalTransistorNmos: 2.78551e+07 muA
** NormalTransistorNmos: 1.00363e+08 muA
** NormalTransistorPmos: -1.7258e+08 muA
** NormalTransistorPmos: -7.48299e+07 muA
** NormalTransistorPmos: -7.48299e+07 muA
** DiodeTransistorNmos: 7.48291e+07 muA
** NormalTransistorNmos: 7.48291e+07 muA
** NormalTransistorPmos: -2.50021e+08 muA
** DiodeTransistorPmos: -2.50022e+08 muA
** NormalTransistorPmos: -7.48289e+07 muA
** NormalTransistorPmos: -7.48289e+07 muA
** NormalTransistorNmos: 3.78487e+08 muA
** NormalTransistorPmos: -3.78486e+08 muA
** DiodeTransistorPmos: -3.78487e+08 muA
** DiodeTransistorNmos: 1.72581e+08 muA
** DiodeTransistorPmos: -2.78559e+07 muA
** NormalTransistorPmos: -2.78569e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.00362e+08 muA


** Expected Voltages: 
** ibias: 3.49701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.575001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.29601  V
** outSourceVoltageBiasXXpXX1: 4.14801  V
** outSourceVoltageBiasXXpXX2: 4.24901  V
** outVoltageBiasXXpXX3: 0.438001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.36001  V
** out1: 0.555001  V
** sourceGCC1: 2.92501  V
** sourceGCC2: 2.92401  V
** inner: 4.14801  V
** inner: 4.24801  V


.END