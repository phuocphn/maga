** Name: two_stage_single_output_op_amp_54_10

.MACRO two_stage_single_output_op_amp_54_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=16e-6
mMainBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=104e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=60e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=21e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=21e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=38e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=38e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=22e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=391e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=60e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
mMainBias14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=141e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=196e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=196e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=496e-6
mMainBias19 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=410e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=503e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=141e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_54_10

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 2.54001 mW
** Area: 13265 (mu_m)^2
** Transit frequency: 3.77001 MHz
** Transit frequency with error factor: 3.77043 MHz
** Slew rate: 4.01151 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 4.46001 V
** VoutMin: 0.210001 V
** VcmMax: 5.17001 V
** VcmMin: 0.790001 V


** Expected Currents: 
** NormalTransistorNmos: 1.35361e+07 muA
** NormalTransistorNmos: 1.52631e+07 muA
** NormalTransistorPmos: -6.02709e+07 muA
** NormalTransistorPmos: -1.90879e+07 muA
** NormalTransistorPmos: -2.89649e+07 muA
** NormalTransistorPmos: -1.90879e+07 muA
** NormalTransistorPmos: -2.89649e+07 muA
** NormalTransistorNmos: 1.90871e+07 muA
** NormalTransistorNmos: 1.90861e+07 muA
** NormalTransistorNmos: 1.90871e+07 muA
** NormalTransistorNmos: 1.90861e+07 muA
** NormalTransistorNmos: 1.97521e+07 muA
** NormalTransistorNmos: 9.87601e+06 muA
** NormalTransistorNmos: 9.87601e+06 muA
** NormalTransistorNmos: 3.51047e+08 muA
** NormalTransistorPmos: -3.51046e+08 muA
** NormalTransistorPmos: -3.51047e+08 muA
** DiodeTransistorNmos: 6.02701e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.35369e+07 muA
** DiodeTransistorPmos: -1.52639e+07 muA


** Expected Voltages: 
** ibias: 0.612001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.04101  V
** out: 2.5  V
** outFirstStage: 4.23601  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.19601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.658001  V
** innerTransistorStack1Load2: 0.452001  V
** innerTransistorStack2Load2: 0.453001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.91901  V
** innerTransconductance: 4.59101  V


.END