** Name: symmetrical_op_amp13

.MACRO symmetrical_op_amp13 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=25e-6
mSecondStage1StageBias5 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mSecondStage1Transconductor6 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor7 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor9 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=111e-6
mMainBias11 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=3e-6 W=301e-6
mSymmetricalFirstStageTransconductor12 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=54e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias13 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mSecondStage1StageBias14 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=1e-6 W=92e-6
mSymmetricalFirstStageTransconductor15 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=54e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp13

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 1.31001 mW
** Area: 1765 (mu_m)^2
** Transit frequency: 3.91001 MHz
** Transit frequency with error factor: 3.91011 MHz
** Slew rate: 3.71473 V/mu_s
** Phase margin: 87.6626°
** CMRR: 153 dB
** negPSRR: 53 dB
** posPSRR: 66 dB
** VoutMax: 3.56001 V
** VoutMin: 0.380001 V
** VcmMax: 4.02001 V
** VcmMin: 0.0100001 V


** Expected Currents: 
** NormalTransistorPmos: -1.22427e+08 muA
** DiodeTransistorNmos: 2.25721e+07 muA
** DiodeTransistorNmos: 2.25721e+07 muA
** NormalTransistorPmos: -4.51469e+07 muA
** NormalTransistorPmos: -2.25729e+07 muA
** NormalTransistorPmos: -2.25729e+07 muA
** NormalTransistorNmos: 3.71921e+07 muA
** NormalTransistorNmos: 3.71931e+07 muA
** NormalTransistorPmos: -3.71929e+07 muA
** DiodeTransistorPmos: -3.71939e+07 muA
** NormalTransistorPmos: -3.71949e+07 muA
** NormalTransistorNmos: 3.71941e+07 muA
** NormalTransistorNmos: 3.71931e+07 muA
** DiodeTransistorNmos: 1.22428e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17601  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.786001  V
** inSourceTransconductanceComplementarySecondStage: 0.577001  V
** inStageBiasComplementarySecondStage: 3.71201  V
** innerComplementarySecondStage: 2.99701  V
** out: 2.5  V
** outFirstStage: 0.577001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21701  V
** innerTransconductance: 0.172001  V
** inner: 0.172001  V


.END