** Name: two_stage_single_output_op_amp_103_2

.MACRO two_stage_single_output_op_amp_103_2 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=150e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=30e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=18e-6
mMainBias6 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=150e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=212e-6
mMainBias9 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=72e-6
mMainBias10 inputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor11 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=106e-6
mTelescopicFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=15e-6
mTelescopicFirstStageStageBias13 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad14 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageTransconductor15 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=353e-6
mTelescopicFirstStageTransconductor16 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=353e-6
mMainBias17 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=513e-6
mSecondStage1StageBias18 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=596e-6
mTelescopicFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=10e-6
mMainBias20 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=90e-6
mTelescopicFirstStageStageBias21 sourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=3e-6 W=189e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11e-12
.EOM two_stage_single_output_op_amp_103_2

** Expected Performance Values: 
** Gain: 146 dB
** Power consumption: 3.25201 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 3.88201 MHz
** Transit frequency with error factor: 3.88207 MHz
** Slew rate: 6.50137 V/mu_s
** Phase margin: 60.1606°
** CMRR: 135 dB
** VoutMax: 4.81001 V
** VoutMin: 0.300001 V
** VcmMax: 3.04001 V
** VcmMin: 0.540001 V


** Expected Currents: 
** NormalTransistorNmos: 1.4666e+08 muA
** NormalTransistorNmos: 2.01361e+07 muA
** NormalTransistorPmos: -3.05699e+07 muA
** NormalTransistorPmos: -1.73491e+08 muA
** NormalTransistorPmos: -2.85709e+07 muA
** NormalTransistorPmos: -2.85709e+07 muA
** DiodeTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorPmos: -2.03804e+08 muA
** NormalTransistorPmos: -2.03803e+08 muA
** NormalTransistorPmos: -2.85719e+07 muA
** NormalTransistorPmos: -2.85719e+07 muA
** NormalTransistorNmos: 2.02445e+08 muA
** NormalTransistorNmos: 2.02444e+08 muA
** NormalTransistorPmos: -2.02444e+08 muA
** DiodeTransistorNmos: 3.05691e+07 muA
** DiodeTransistorNmos: 1.73492e+08 muA
** DiodeTransistorPmos: -1.46659e+08 muA
** DiodeTransistorPmos: -2.01369e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXpXX1: 2.04101  V
** inputVoltageBiasXXpXX2: 3.51301  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.560001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.27701  V
** innerStageBias: 4.50101  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.00601  V
** sourceGCC2: 3.00301  V
** innerTransconductance: 0.150001  V


.END