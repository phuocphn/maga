** Name: two_stage_single_output_op_amp_51_3

.MACRO two_stage_single_output_op_amp_51_3 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=94e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=31e-6
mMainBias3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=46e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=47e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=94e-6
mFoldedCascodeFirstStageTransconductor6 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=32e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=32e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=8e-6 W=116e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=263e-6
mFoldedCascodeFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=5e-6 W=43e-6
mMainBias11 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=241e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 outInputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=6e-6 W=21e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=27e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=27e-6
mSecondStage1StageBias15 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=482e-6
mSecondStage1StageBias16 out outInputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=6e-6 W=595e-6
mFoldedCascodeFirstStageLoad17 outFirstStage outInputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=6e-6 W=21e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.70001e-12
.EOM two_stage_single_output_op_amp_51_3

** Expected Performance Values: 
** Gain: 118 dB
** Power consumption: 4.86801 mW
** Area: 14783 (mu_m)^2
** Transit frequency: 3.99601 MHz
** Transit frequency with error factor: 3.99581 MHz
** Slew rate: 3.8319 V/mu_s
** Phase margin: 60.1606°
** CMRR: 130 dB
** VoutMax: 3.02001 V
** VoutMin: 0.540001 V
** VcmMax: 4.66001 V
** VcmMin: 0.800001 V


** Expected Currents: 
** NormalTransistorNmos: 7.78411e+07 muA
** NormalTransistorPmos: -2.57549e+07 muA
** NormalTransistorPmos: -4.41529e+07 muA
** NormalTransistorPmos: -2.57539e+07 muA
** NormalTransistorPmos: -4.41519e+07 muA
** NormalTransistorNmos: 2.57541e+07 muA
** NormalTransistorNmos: 2.57531e+07 muA
** DiodeTransistorNmos: 2.57541e+07 muA
** NormalTransistorNmos: 3.67941e+07 muA
** NormalTransistorNmos: 1.83971e+07 muA
** NormalTransistorNmos: 1.83971e+07 muA
** NormalTransistorNmos: 7.97511e+08 muA
** NormalTransistorPmos: -7.9751e+08 muA
** NormalTransistorPmos: -7.97511e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.78419e+07 muA
** DiodeTransistorPmos: -7.78429e+07 muA


** Expected Voltages: 
** ibias: 0.579001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.943001  V
** outInputVoltageBiasXXpXX1: 2.37801  V
** outSourceVoltageBiasXXpXX1: 3.69201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** out1: 1.14801  V
** sourceGCC1: 3.58101  V
** sourceGCC2: 3.58101  V
** sourceTransconductance: 1.87601  V
** innerStageBias: 3.61001  V


.END