** Name: two_stage_single_output_op_amp_44_8

.MACRO two_stage_single_output_op_amp_44_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=126e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=126e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=105e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=56e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=97e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=97e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=516e-6
mFoldedCascodeFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=56e-6
mFoldedCascodeFirstStageLoad11 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=105e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=135e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=135e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=229e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=443e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=401e-6
mFoldedCascodeFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=124e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9e-12
.EOM two_stage_single_output_op_amp_44_8

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 4.51001 mW
** Area: 10282 (mu_m)^2
** Transit frequency: 3.43001 MHz
** Transit frequency with error factor: 3.42961 MHz
** Slew rate: 6.72479 V/mu_s
** Phase margin: 60.1606°
** CMRR: 141 dB
** VoutMax: 4.43001 V
** VoutMin: 0.720001 V
** VcmMax: 3.87001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.19992e+08 muA
** NormalTransistorNmos: 6.08521e+07 muA
** NormalTransistorNmos: 9.23751e+07 muA
** NormalTransistorNmos: 6.08511e+07 muA
** NormalTransistorNmos: 9.23751e+07 muA
** NormalTransistorPmos: -6.08529e+07 muA
** NormalTransistorPmos: -6.08519e+07 muA
** DiodeTransistorPmos: -6.08529e+07 muA
** NormalTransistorPmos: -6.30459e+07 muA
** NormalTransistorPmos: -3.15229e+07 muA
** NormalTransistorPmos: -3.15229e+07 muA
** NormalTransistorNmos: 5.77161e+08 muA
** NormalTransistorNmos: 5.7716e+08 muA
** NormalTransistorPmos: -5.7716e+08 muA
** DiodeTransistorNmos: 1.19993e+08 muA
** DiodeTransistorNmos: 1.19993e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11001  V
** out: 2.5  V
** outFirstStage: 3.86601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.25601  V
** out1: 3.52601  V
** sourceGCC1: 0.544001  V
** sourceGCC2: 0.544001  V
** sourceTransconductance: 3.38601  V
** innerStageBias: 0.542001  V


.END