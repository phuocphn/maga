** Name: two_stage_single_output_op_amp_45_6

.MACRO two_stage_single_output_op_amp_45_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=22e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=51e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
mMainBias5 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=12e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=12e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=197e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=27e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=79e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=79e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=279e-6
mMainBias12 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=22e-6
mMainBias13 inputVoltageBiasXXpXX3 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=11e-6
mSecondStage1Transconductor14 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=259e-6
mFoldedCascodeFirstStageLoad15 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=27e-6
mMainBias16 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=17e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=51e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=17e-6
mFoldedCascodeFirstStageStageBias20 FirstStageYsourceTransconductance inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=72e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=12e-6
mMainBias22 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=377e-6
mSecondStage1StageBias23 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=197e-6
mFoldedCascodeFirstStageLoad24 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=8e-6 W=334e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_45_6

** Expected Performance Values: 
** Gain: 174 dB
** Power consumption: 1.91901 mW
** Area: 14887 (mu_m)^2
** Transit frequency: 2.63801 MHz
** Transit frequency with error factor: 2.63808 MHz
** Slew rate: 4.4324 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 3.44001 V
** VoutMin: 0.340001 V
** VcmMax: 3.63001 V
** VcmMin: -0.359999 V


** Expected Currents: 
** NormalTransistorNmos: 7.63201e+06 muA
** NormalTransistorNmos: 1.00751e+07 muA
** NormalTransistorNmos: 5.00501e+06 muA
** NormalTransistorPmos: -1.56825e+08 muA
** NormalTransistorNmos: 2.06871e+07 muA
** NormalTransistorNmos: 3.54641e+07 muA
** NormalTransistorNmos: 2.06871e+07 muA
** NormalTransistorNmos: 3.54641e+07 muA
** DiodeTransistorPmos: -2.06879e+07 muA
** NormalTransistorPmos: -2.06879e+07 muA
** NormalTransistorPmos: -2.06879e+07 muA
** NormalTransistorPmos: -2.95529e+07 muA
** NormalTransistorPmos: -1.47759e+07 muA
** NormalTransistorPmos: -1.47759e+07 muA
** NormalTransistorNmos: 1.23326e+08 muA
** NormalTransistorNmos: 1.23325e+08 muA
** NormalTransistorPmos: -1.23325e+08 muA
** DiodeTransistorPmos: -1.23326e+08 muA
** DiodeTransistorNmos: 1.56826e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.63299e+06 muA
** NormalTransistorPmos: -7.63399e+06 muA
** DiodeTransistorPmos: -1.00759e+07 muA
** DiodeTransistorPmos: -5.00599e+06 muA


** Expected Voltages: 
** ibias: 0.612001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.00201  V
** inputVoltageBiasXXpXX2: 3.68601  V
** inputVoltageBiasXXpXX3: 4.00601  V
** out: 2.5  V
** outFirstStage: 0.597001  V
** outInputVoltageBiasXXpXX1: 2.87801  V
** outSourceVoltageBiasXXpXX1: 3.93901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.41601  V
** out1: 4.17401  V
** sourceGCC1: 0.407001  V
** sourceGCC2: 0.407001  V
** sourceTransconductance: 3.44501  V
** innerTransconductance: 0.447001  V
** inner: 3.93901  V


.END