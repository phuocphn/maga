** Name: two_stage_single_output_op_amp_198_11

.MACRO two_stage_single_output_op_amp_198_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=1e-6 W=14e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=15e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=89e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=121e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=16e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=71e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=121e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=89e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=303e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=14e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=71e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=355e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=21e-6
mSimpleFirstStageLoad19 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=571e-6
mSimpleFirstStageLoad20 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=571e-6
mSimpleFirstStageLoad21 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=204e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSecondStage1Transconductor23 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=598e-6
mSimpleFirstStageLoad24 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=204e-6
mMainBias25 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=38e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.80001e-12
.EOM two_stage_single_output_op_amp_198_11

** Expected Performance Values: 
** Gain: 150 dB
** Power consumption: 8.38901 mW
** Area: 13824 (mu_m)^2
** Transit frequency: 8.13101 MHz
** Transit frequency with error factor: 8.12532 MHz
** Slew rate: 7.66371 V/mu_s
** Phase margin: 60.1606°
** CMRR: 121 dB
** VoutMax: 4.62001 V
** VoutMin: 0.770001 V
** VcmMax: 4.66001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 2.33528e+08 muA
** NormalTransistorNmos: 1.40111e+07 muA
** NormalTransistorPmos: -3.35379e+07 muA
** DiodeTransistorNmos: 4.73132e+08 muA
** DiodeTransistorNmos: 4.73131e+08 muA
** NormalTransistorNmos: 4.7313e+08 muA
** NormalTransistorNmos: 4.73131e+08 muA
** NormalTransistorPmos: -4.9567e+08 muA
** NormalTransistorPmos: -4.95669e+08 muA
** NormalTransistorPmos: -4.95668e+08 muA
** NormalTransistorPmos: -4.95669e+08 muA
** NormalTransistorNmos: 4.50771e+07 muA
** DiodeTransistorNmos: 4.50761e+07 muA
** NormalTransistorNmos: 2.25391e+07 muA
** NormalTransistorNmos: 2.25391e+07 muA
** NormalTransistorNmos: 3.95348e+08 muA
** NormalTransistorNmos: 3.95347e+08 muA
** NormalTransistorPmos: -3.95347e+08 muA
** NormalTransistorPmos: -3.95348e+08 muA
** DiodeTransistorNmos: 3.35371e+07 muA
** NormalTransistorNmos: 3.35361e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.33527e+08 muA
** DiodeTransistorPmos: -1.40119e+07 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.24401  V
** outInputVoltageBiasXXnXX1: 1.20901  V
** outSourceVoltageBiasXXnXX1: 0.605001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.05301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack1Load2: 4.61701  V
** innerTransistorStack2Load1: 1.15601  V
** innerTransistorStack2Load2: 4.61701  V
** out1: 2.19501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.495001  V
** innerTransconductance: 4.44201  V
** inner: 0.603001  V


.END