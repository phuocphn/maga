** Name: two_stage_single_output_op_amp_144_7

.MACRO two_stage_single_output_op_amp_144_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=91e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=438e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=28e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
mMainBias8 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=199e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=560e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=6e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=28e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=95e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=95e-6
mSimpleFirstStageLoad14 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=17e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=387e-6
mSimpleFirstStageLoad16 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=17e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_144_7

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 4.28301 mW
** Area: 7238 (mu_m)^2
** Transit frequency: 3.21701 MHz
** Transit frequency with error factor: 3.21434 MHz
** Slew rate: 3.50059 V/mu_s
** Phase margin: 61.3065°
** CMRR: 108 dB
** VoutMax: 4.25 V
** VoutMin: 0.190001 V
** VcmMax: 4.65001 V
** VcmMin: 0.770001 V


** Expected Currents: 
** NormalTransistorNmos: 2.00122e+08 muA
** NormalTransistorNmos: 3.46521e+07 muA
** NormalTransistorNmos: 3.46511e+07 muA
** DiodeTransistorNmos: 3.46521e+07 muA
** NormalTransistorPmos: -4.25519e+07 muA
** NormalTransistorPmos: -4.25519e+07 muA
** NormalTransistorPmos: -4.25509e+07 muA
** NormalTransistorPmos: -4.25519e+07 muA
** NormalTransistorNmos: 1.57991e+07 muA
** NormalTransistorNmos: 7.89901e+06 muA
** NormalTransistorNmos: 7.89901e+06 muA
** NormalTransistorNmos: 5.61338e+08 muA
** NormalTransistorPmos: -5.61337e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.00121e+08 muA
** DiodeTransistorPmos: -2.00122e+08 muA


** Expected Voltages: 
** ibias: 0.593001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.14901  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.21101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.04801  V
** innerTransistorStack1Load2: 4.24001  V
** innerTransistorStack2Load2: 4.24001  V
** out1: 2.09501  V
** sourceTransconductance: 1.92101  V


.END