** Name: two_stage_single_output_op_amp_62_6

.MACRO two_stage_single_output_op_amp_62_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=7e-6 W=60e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=13e-6
mMainBias5 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=5e-6 W=28e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=53e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=473e-6
mMainBias8 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=17e-6
mMainBias9 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=9e-6 W=26e-6
mFoldedCascodeFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=32e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=39e-6
mFoldedCascodeFirstStageLoad12 FirstStageYsourceGCC2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=39e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=412e-6
mSecondStage1Transconductor14 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=186e-6
mFoldedCascodeFirstStageLoad15 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=32e-6
mMainBias16 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mMainBias17 outInputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=19e-6
mMainBias18 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mMainBias19 outVoltageBiasXXpXX3 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=35e-6
mFoldedCascodeFirstStageLoad20 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=7e-6 W=60e-6
mFoldedCascodeFirstStageTransconductor21 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=78e-6
mFoldedCascodeFirstStageTransconductor22 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=78e-6
mFoldedCascodeFirstStageStageBias23 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=53e-6
mMainBias24 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=13e-6
mMainBias25 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=28e-6
mSecondStage1StageBias26 out outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=5e-6 W=473e-6
mFoldedCascodeFirstStageLoad27 outFirstStage outVoltageBiasXXpXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=9e-6 W=283e-6
mMainBias28 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=208e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.20001e-12
.EOM two_stage_single_output_op_amp_62_6

** Expected Performance Values: 
** Gain: 178 dB
** Power consumption: 2.34101 mW
** Area: 14987 (mu_m)^2
** Transit frequency: 3.69101 MHz
** Transit frequency with error factor: 3.69078 MHz
** Slew rate: 3.55223 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 3.64001 V
** VoutMin: 0.510001 V
** VcmMax: 3.07001 V
** VcmMin: -0.369999 V


** Expected Currents: 
** NormalTransistorNmos: 5.75101e+06 muA
** NormalTransistorNmos: 6.57201e+06 muA
** NormalTransistorNmos: 1.56931e+07 muA
** NormalTransistorNmos: 2.93311e+07 muA
** NormalTransistorPmos: -7.15e+07 muA
** NormalTransistorNmos: 1.86881e+07 muA
** NormalTransistorNmos: 3.20371e+07 muA
** NormalTransistorNmos: 1.86881e+07 muA
** NormalTransistorNmos: 3.20371e+07 muA
** DiodeTransistorPmos: -1.86889e+07 muA
** NormalTransistorPmos: -1.86889e+07 muA
** NormalTransistorPmos: -1.86889e+07 muA
** NormalTransistorPmos: -2.66969e+07 muA
** DiodeTransistorPmos: -2.66979e+07 muA
** NormalTransistorPmos: -1.33479e+07 muA
** NormalTransistorPmos: -1.33479e+07 muA
** NormalTransistorNmos: 2.65305e+08 muA
** NormalTransistorNmos: 2.65306e+08 muA
** NormalTransistorPmos: -2.65304e+08 muA
** DiodeTransistorPmos: -2.65305e+08 muA
** DiodeTransistorNmos: 7.14991e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.75199e+06 muA
** DiodeTransistorPmos: -6.57299e+06 muA
** NormalTransistorPmos: -6.57399e+06 muA
** DiodeTransistorPmos: -1.56939e+07 muA
** NormalTransistorPmos: -1.56949e+07 muA
** DiodeTransistorPmos: -2.93319e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.601001  V
** outInputVoltageBiasXXpXX1: 3.28801  V
** outInputVoltageBiasXXpXX2: 3.07601  V
** outSourceVoltageBiasXXpXX1: 4.14401  V
** outSourceVoltageBiasXXpXX2: 4.03801  V
** outVoltageBiasXXnXX1: 1.00601  V
** outVoltageBiasXXpXX0: 4.16001  V
** outVoltageBiasXXpXX3: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.43201  V
** out1: 4.08501  V
** sourceGCC1: 0.398001  V
** sourceGCC2: 0.398001  V
** sourceTransconductance: 3.28201  V
** innerTransconductance: 0.282001  V
** inner: 4.14201  V
** inner: 4.03501  V


.END