** Name: two_stage_single_output_op_amp_47_5

.MACRO two_stage_single_output_op_amp_47_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=16e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mMainBias3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mMainBias4 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=10e-6 W=78e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=6e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=307e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
mMainBias10 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=106e-6
mMainBias11 inputVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=37e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=172e-6
mFoldedCascodeFirstStageLoad13 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=26e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=24e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=19e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=29e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=152e-6
mFoldedCascodeFirstStageTransconductor19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=152e-6
mFoldedCascodeFirstStageStageBias20 FirstStageYsourceTransconductance inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=10e-6 W=119e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=307e-6
mFoldedCascodeFirstStageLoad23 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=19e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.30001e-12
.EOM two_stage_single_output_op_amp_47_5

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 3.03801 mW
** Area: 12295 (mu_m)^2
** Transit frequency: 3.40701 MHz
** Transit frequency with error factor: 3.40665 MHz
** Slew rate: 3.934 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 3 V
** VoutMin: 0.540001 V
** VcmMax: 3.93001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 9.17101e+06 muA
** NormalTransistorNmos: 4.06121e+07 muA
** NormalTransistorNmos: 1.40951e+07 muA
** NormalTransistorNmos: 2.09031e+07 muA
** NormalTransistorNmos: 3.16171e+07 muA
** NormalTransistorNmos: 2.09031e+07 muA
** NormalTransistorNmos: 3.16171e+07 muA
** NormalTransistorPmos: -2.09039e+07 muA
** NormalTransistorPmos: -2.09049e+07 muA
** NormalTransistorPmos: -2.09039e+07 muA
** NormalTransistorPmos: -2.09049e+07 muA
** NormalTransistorPmos: -2.14309e+07 muA
** NormalTransistorPmos: -1.07149e+07 muA
** NormalTransistorPmos: -1.07149e+07 muA
** NormalTransistorNmos: 4.70534e+08 muA
** NormalTransistorPmos: -4.70533e+08 muA
** DiodeTransistorPmos: -4.70534e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.17199e+06 muA
** NormalTransistorPmos: -9.17299e+06 muA
** DiodeTransistorPmos: -4.06129e+07 muA
** DiodeTransistorPmos: -1.40959e+07 muA


** Expected Voltages: 
** ibias: 1.15201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.68601  V
** inputVoltageBiasXXpXX3: 4.11701  V
** out: 2.5  V
** outFirstStage: 0.947001  V
** outInputVoltageBiasXXpXX1: 2.43601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.71601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.23601  V
** innerTransistorStack1Load2: 4.60001  V
** innerTransistorStack2Load2: 4.60001  V
** sourceGCC1: 0.528001  V
** sourceGCC2: 0.528001  V
** sourceTransconductance: 3.25201  V
** inner: 3.71301  V


.END