** Design view name: schematic
.GLOBAL vdd! gnd!

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: CascodeSymmetricalCMOSOTA
** Cell name: cascodeSymmetricalCMOSOTA
** View name: schematic
c1 outFirstStage out 
c2 outSecondStage out 
m1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 gnd! gnd! nmos
m2 outInputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 gnd! gnd! nmos
m3 outVoltageBiasXXnXX0 ibias vdd! vdd! pmos
m4 inputVoltageBiasXXnXX1 ibias vdd! vdd! pmos
m5 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m6 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 gnd! gnd! nmos
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 gnd! gnd! nmos
m9 FirstStageYsourceTransconductance ibias vdd! vdd! pmos
m10 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out gnd! 
m12 outSecondStage outFirstStage gnd! gnd! nmos
m13 outSecondStage outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m14 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 vdd! vdd! pmos
m15 out outSecondStage gnd! gnd! nmos
m16 out outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m17 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 vdd! vdd! pmos
m18 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 gnd! gnd! nmos
m19 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 gnd! gnd! nmos
m20 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 vdd! vdd! pmos
m22 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m23 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 vdd! vdd! pmos
m24 ibias ibias vdd! vdd! pmos
.END