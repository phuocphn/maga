** Name: two_stage_single_output_op_amp_89_7

.MACRO two_stage_single_output_op_amp_89_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=11e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=89e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=8e-6
mTelescopicFirstStageLoad5 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=7e-6 W=78e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=89e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=89e-6
mSecondStage1StageBias8 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=78e-6
mMainBias10 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mTelescopicFirstStageLoad11 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=55e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=83e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=83e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=105e-6
mMainBias15 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=405e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=179e-6
mTelescopicFirstStageLoad17 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=55e-6
mTelescopicFirstStageStageBias18 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=490e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.8001e-12
.EOM two_stage_single_output_op_amp_89_7

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 8.87701 mW
** Area: 12000 (mu_m)^2
** Transit frequency: 2.75501 MHz
** Transit frequency with error factor: 2.75524 MHz
** Slew rate: 4.73636 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 3.39001 V
** VoutMin: 0.25 V
** VcmMax: 4.03001 V
** VcmMin: -0.209999 V


** Expected Currents: 
** NormalTransistorNmos: 1.36031e+07 muA
** NormalTransistorPmos: -1.18549e+07 muA
** NormalTransistorPmos: -4.56019e+07 muA
** NormalTransistorPmos: -2.12239e+07 muA
** NormalTransistorPmos: -2.12239e+07 muA
** NormalTransistorNmos: 2.12231e+07 muA
** NormalTransistorNmos: 2.12221e+07 muA
** NormalTransistorNmos: 2.12231e+07 muA
** NormalTransistorNmos: 2.12221e+07 muA
** NormalTransistorPmos: -5.60529e+07 muA
** NormalTransistorPmos: -2.12249e+07 muA
** NormalTransistorPmos: -2.12249e+07 muA
** NormalTransistorNmos: 1.64193e+09 muA
** NormalTransistorPmos: -1.64192e+09 muA
** DiodeTransistorNmos: 1.18541e+07 muA
** DiodeTransistorNmos: 4.56011e+07 muA
** DiodeTransistorPmos: -1.36039e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXnXX2: 0.658001  V
** out: 2.5  V
** outFirstStage: 2.82601  V
** outVoltageBiasXXpXX1: 2.26901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.27101  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 3.04001  V
** sourceGCC2: 3.04001  V


.END