** Name: symmetrical_op_amp154

.MACRO symmetrical_op_amp154 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=12e-6
mMainBias2 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=20e-6
mSecondStage1StageBias3 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=38e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=3e-6 W=38e-6
mSymmetricalFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=110e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=44e-6
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=44e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=122e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=122e-6
mSymmetricalFirstStageLoad10 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=38e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=8e-6 W=82e-6
mSecondStage1Transconductor12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=8e-6 W=82e-6
mSymmetricalFirstStageLoad13 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=8e-6 W=38e-6
mSymmetricalFirstStageStageBias14 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=110e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias15 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=38e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mSymmetricalFirstStageTransconductor17 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=99e-6
mSecondStage1StageBias18 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=3e-6 W=38e-6
mSymmetricalFirstStageTransconductor19 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=99e-6
mMainBias20 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp154

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 1.28201 mW
** Area: 5388 (mu_m)^2
** Transit frequency: 4.38801 MHz
** Transit frequency with error factor: 4.38828 MHz
** Slew rate: 7.73494 V/mu_s
** Phase margin: 65.8902°
** CMRR: 140 dB
** negPSRR: 43 dB
** posPSRR: 60 dB
** VoutMax: 3.26001 V
** VoutMin: 0.450001 V
** VcmMax: 3.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.54749e+07 muA
** NormalTransistorNmos: 2.80231e+07 muA
** NormalTransistorNmos: 2.80221e+07 muA
** NormalTransistorNmos: 2.80231e+07 muA
** NormalTransistorNmos: 2.80221e+07 muA
** NormalTransistorPmos: -5.60469e+07 muA
** DiodeTransistorPmos: -5.60459e+07 muA
** NormalTransistorPmos: -2.80239e+07 muA
** NormalTransistorPmos: -2.80239e+07 muA
** NormalTransistorNmos: 7.74541e+07 muA
** NormalTransistorNmos: 7.74551e+07 muA
** NormalTransistorPmos: -7.74549e+07 muA
** DiodeTransistorPmos: -7.74559e+07 muA
** DiodeTransistorPmos: -7.74549e+07 muA
** NormalTransistorPmos: -7.74559e+07 muA
** NormalTransistorNmos: 7.74541e+07 muA
** NormalTransistorNmos: 7.74551e+07 muA
** DiodeTransistorNmos: 2.54741e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.28801  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 3.84901  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 2.69801  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.853001  V
** outSourceVoltageBiasXXpXX1: 4.14501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.183001  V
** innerTransistorStack2Load1: 0.183001  V
** sourceTransconductance: 3.34501  V
** innerTransconductance: 0.150001  V
** inner: 3.84501  V
** inner: 0.150001  V
** inner: 4.14101  V


.END