** Name: two_stage_single_output_op_amp_106_3

.MACRO two_stage_single_output_op_amp_106_3 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=64e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=64e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=280e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos4 L=4e-6 W=17e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=154e-6
mMainBias7 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=10e-6
mTelescopicFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=64e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=415e-6
mTelescopicFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=64e-6
mMainBias12 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=21e-6
mMainBias13 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=186e-6
mTelescopicFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=9e-6
mTelescopicFirstStageTransconductor15 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=36e-6
mTelescopicFirstStageTransconductor16 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=36e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=4e-6 W=138e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias19 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=4e-6 W=21e-6
mSecondStage1StageBias20 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=4e-6 W=599e-6
mTelescopicFirstStageLoad21 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=9e-6
mTelescopicFirstStageStageBias22 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=154e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_106_3

** Expected Performance Values: 
** Gain: 133 dB
** Power consumption: 2.45701 mW
** Area: 14909 (mu_m)^2
** Transit frequency: 2.93201 MHz
** Transit frequency with error factor: 2.93242 MHz
** Slew rate: 13.8482 V/mu_s
** Phase margin: 65.8902°
** CMRR: 130 dB
** VoutMax: 3.32001 V
** VoutMin: 0.300001 V
** VcmMax: 3.25 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorNmos: 4.03301e+06 muA
** NormalTransistorNmos: 3.56611e+07 muA
** NormalTransistorPmos: -5.34469e+07 muA
** NormalTransistorPmos: -1.35459e+07 muA
** NormalTransistorPmos: -1.35459e+07 muA
** DiodeTransistorNmos: 1.35451e+07 muA
** DiodeTransistorNmos: 1.35451e+07 muA
** NormalTransistorNmos: 1.35451e+07 muA
** NormalTransistorNmos: 1.35451e+07 muA
** NormalTransistorPmos: -6.27569e+07 muA
** DiodeTransistorPmos: -6.27579e+07 muA
** NormalTransistorPmos: -1.35469e+07 muA
** NormalTransistorPmos: -1.35469e+07 muA
** NormalTransistorNmos: 3.51228e+08 muA
** NormalTransistorPmos: -3.51227e+08 muA
** NormalTransistorPmos: -3.51226e+08 muA
** DiodeTransistorNmos: 5.34461e+07 muA
** DiodeTransistorPmos: -4.03399e+06 muA
** NormalTransistorPmos: -4.03499e+06 muA
** DiodeTransistorPmos: -3.56619e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.75701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outInputVoltageBiasXXpXX1: 3.57001  V
** outSourceVoltageBiasXXpXX1: 4.28501  V
** outSourceVoltageBiasXXpXX3: 3.68501  V
** outVoltageBiasXXpXX2: 1.64701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.38701  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 2.98201  V
** sourceGCC2: 2.97501  V
** innerStageBias: 3.68201  V
** inner: 4.28401  V


.END