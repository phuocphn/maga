** Name: two_stage_single_output_op_amp_198_8

.MACRO two_stage_single_output_op_amp_198_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=9e-6 W=17e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=27e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=253e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=22e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=8e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=20e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=464e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=253e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=316e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=9e-6 W=17e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=20e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=47e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=47e-6
mSimpleFirstStageLoad19 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=314e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=44e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=388e-6
mSimpleFirstStageLoad22 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=314e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=391e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.20001e-12
.EOM two_stage_single_output_op_amp_198_8

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 9.98401 mW
** Area: 6672 (mu_m)^2
** Transit frequency: 4.26801 MHz
** Transit frequency with error factor: 4.26662 MHz
** Slew rate: 4.02264 V/mu_s
** Phase margin: 60.1606°
** CMRR: 110 dB
** VoutMax: 4.25 V
** VoutMin: 0.810001 V
** VcmMax: 4.77001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorPmos: -4.89906e+08 muA
** NormalTransistorPmos: -5.55239e+07 muA
** DiodeTransistorNmos: 4.63921e+07 muA
** DiodeTransistorNmos: 4.63931e+07 muA
** NormalTransistorNmos: 4.63921e+07 muA
** NormalTransistorNmos: 4.63931e+07 muA
** NormalTransistorPmos: -5.90909e+07 muA
** NormalTransistorPmos: -5.90919e+07 muA
** NormalTransistorPmos: -5.90909e+07 muA
** NormalTransistorPmos: -5.90919e+07 muA
** NormalTransistorNmos: 2.53951e+07 muA
** DiodeTransistorNmos: 2.53941e+07 muA
** NormalTransistorNmos: 1.26981e+07 muA
** NormalTransistorNmos: 1.26981e+07 muA
** NormalTransistorNmos: 1.31318e+09 muA
** NormalTransistorNmos: 1.31318e+09 muA
** NormalTransistorPmos: -1.31317e+09 muA
** DiodeTransistorNmos: 4.89907e+08 muA
** NormalTransistorNmos: 4.89908e+08 muA
** DiodeTransistorNmos: 5.55231e+07 muA
** DiodeTransistorNmos: 5.55241e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.14801  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.11401  V
** outSourceVoltageBiasXXnXX1: 0.557001  V
** outSourceVoltageBiasXXnXX2: 0.587001  V
** outSourceVoltageBiasXXpXX1: 3.97601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.14901  V
** innerTransistorStack1Load2: 3.87601  V
** innerTransistorStack2Load1: 1.14901  V
** innerTransistorStack2Load2: 3.87601  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.521001  V
** inner: 0.558001  V


.END