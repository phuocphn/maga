** Name: two_stage_single_output_op_amp_196_9

.MACRO two_stage_single_output_op_amp_196_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=11e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=15e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=6e-6
mMainBias4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=4e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=143e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=331e-6
mMainBias7 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=11e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=28e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=143e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=331e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=15e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=28e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=304e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=532e-6
mSimpleFirstStageLoad18 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=304e-6
mMainBias19 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias20 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=69e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.3001e-12
.EOM two_stage_single_output_op_amp_196_9

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 14.9991 mW
** Area: 6609 (mu_m)^2
** Transit frequency: 5.83901 MHz
** Transit frequency with error factor: 5.82983 MHz
** Slew rate: 5.50283 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 1.63001 V
** VcmMax: 5.25 V
** VcmMin: 1.42001 V


** Expected Currents: 
** NormalTransistorPmos: -4.52999e+06 muA
** NormalTransistorPmos: -3.16779e+07 muA
** DiodeTransistorNmos: 8.55561e+07 muA
** DiodeTransistorNmos: 8.55551e+07 muA
** NormalTransistorNmos: 8.55541e+07 muA
** NormalTransistorNmos: 8.55551e+07 muA
** NormalTransistorPmos: -1.38884e+08 muA
** NormalTransistorPmos: -1.38884e+08 muA
** NormalTransistorNmos: 1.0666e+08 muA
** DiodeTransistorNmos: 1.06659e+08 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 2.66593e+09 muA
** DiodeTransistorNmos: 2.66593e+09 muA
** NormalTransistorPmos: -2.66592e+09 muA
** DiodeTransistorNmos: 4.52901e+06 muA
** NormalTransistorNmos: 4.52801e+06 muA
** DiodeTransistorNmos: 3.16771e+07 muA
** NormalTransistorNmos: 3.16761e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.27001  V
** outInputVoltageBiasXXnXX2: 2.03801  V
** outSourceVoltageBiasXXnXX1: 0.636001  V
** outSourceVoltageBiasXXnXX2: 1.01901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15101  V
** innerTransistorStack2Load1: 1.15201  V
** out1: 2.19501  V
** sourceTransconductance: 1.94501  V
** inner: 0.633001  V
** inner: 1.01901  V


.END