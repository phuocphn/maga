** Name: two_stage_single_output_op_amp_54_7

.MACRO two_stage_single_output_op_amp_54_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=96e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=66e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=10e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=24e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=105e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=26e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=26e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=406e-6
mFoldedCascodeFirstStageLoad12 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=105e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=145e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=106e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=106e-6
mMainBias16 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=499e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=88e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=145e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=569e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.90001e-12
.EOM two_stage_single_output_op_amp_54_7

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 7.28301 mW
** Area: 6548 (mu_m)^2
** Transit frequency: 3.70301 MHz
** Transit frequency with error factor: 3.70251 MHz
** Slew rate: 3.69634 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 4.25 V
** VoutMin: 0.160001 V
** VcmMax: 5.19001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorPmos: -2.41818e+08 muA
** NormalTransistorPmos: -2.11158e+08 muA
** NormalTransistorPmos: -2.94439e+07 muA
** NormalTransistorPmos: -4.50479e+07 muA
** NormalTransistorPmos: -2.94439e+07 muA
** NormalTransistorPmos: -4.50479e+07 muA
** NormalTransistorNmos: 2.94431e+07 muA
** NormalTransistorNmos: 2.94421e+07 muA
** NormalTransistorNmos: 2.94431e+07 muA
** NormalTransistorNmos: 2.94421e+07 muA
** NormalTransistorNmos: 3.12051e+07 muA
** NormalTransistorNmos: 1.56031e+07 muA
** NormalTransistorNmos: 1.56031e+07 muA
** NormalTransistorNmos: 8.93499e+08 muA
** NormalTransistorPmos: -8.93498e+08 muA
** DiodeTransistorNmos: 2.41819e+08 muA
** DiodeTransistorNmos: 2.11159e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.567001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.21901  V
** outVoltageBiasXXnXX1: 1.02801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.656001  V
** innerTransistorStack1Load2: 0.450001  V
** innerTransistorStack2Load2: 0.451001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.92601  V


.END