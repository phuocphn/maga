** Name: symmetrical_op_amp27

.MACRO symmetrical_op_amp27 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=26e-6
mSecondStage1StageBias2 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mSecondStage1StageBias3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
mSymmetricalFirstStageLoad4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=86e-6
mSymmetricalFirstStageLoad5 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=86e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=6e-6 W=600e-6
mMainBias7 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos4 L=6e-6 W=33e-6
mSymmetricalFirstStageTransconductor8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=180e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias9 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mSecondStage1StageBias10 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos4 L=1e-6 W=13e-6
mSymmetricalFirstStageTransconductor11 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=180e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=125e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor13 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=125e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=4e-6 W=170e-6
mSecondStage1Transconductor15 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=170e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp27

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 2.99601 mW
** Area: 7285 (mu_m)^2
** Transit frequency: 15.375 MHz
** Transit frequency with error factor: 15.3746 MHz
** Slew rate: 17.1554 V/mu_s
** Phase margin: 61.3065°
** CMRR: 141 dB
** negPSRR: 56 dB
** posPSRR: 47 dB
** VoutMax: 4.25 V
** VoutMin: 1.26001 V
** VcmMax: 4.57001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorNmos: 1.26901e+07 muA
** DiodeTransistorPmos: -1.16394e+08 muA
** DiodeTransistorPmos: -1.16394e+08 muA
** NormalTransistorNmos: 2.32788e+08 muA
** NormalTransistorNmos: 1.16395e+08 muA
** NormalTransistorNmos: 1.16395e+08 muA
** NormalTransistorNmos: 1.71877e+08 muA
** DiodeTransistorNmos: 1.71876e+08 muA
** NormalTransistorPmos: -1.71876e+08 muA
** NormalTransistorPmos: -1.71875e+08 muA
** NormalTransistorNmos: 1.71877e+08 muA
** NormalTransistorPmos: -1.71876e+08 muA
** NormalTransistorPmos: -1.71875e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.26909e+07 muA


** Expected Voltages: 
** ibias: 0.570001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 4.16001  V
** inStageBiasComplementarySecondStage: 0.865001  V
** innerComplementarySecondStage: 1.66401  V
** out: 2.5  V
** outFirstStage: 4.16001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.92001  V
** innerTransconductance: 4.72401  V
** inner: 4.72401  V


.END