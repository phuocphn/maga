** Name: symmetrical_op_amp81

.MACRO symmetrical_op_amp81 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=20e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSymmetricalFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mSecondStage1StageBias4 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSymmetricalFirstStageLoad5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=91e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=32e-6
mSymmetricalFirstStageLoad7 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=91e-6
mSymmetricalFirstStageStageBias8 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=600e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=153e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias10 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=153e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=20e-6
mMainBias12 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=20e-6
mSymmetricalFirstStageTransconductor13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=22e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias14 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=2e-6 W=64e-6
mMainBias15 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSecondStage1StageBias16 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=67e-6
mSymmetricalFirstStageTransconductor17 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=22e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=103e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor19 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=103e-6
mMainBias20 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=600e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor21 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=3e-6 W=496e-6
mSecondStage1Transconductor22 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=496e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp81

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 3.48001 mW
** Area: 14680 (mu_m)^2
** Transit frequency: 3.55401 MHz
** Transit frequency with error factor: 3.55443 MHz
** Slew rate: 16.9698 V/mu_s
** Phase margin: 83.0789°
** CMRR: 133 dB
** negPSRR: 55 dB
** posPSRR: 41 dB
** VoutMax: 4.46001 V
** VoutMin: 0.410001 V
** VcmMax: 4.54001 V
** VcmMin: 1.86001 V


** Expected Currents: 
** NormalTransistorNmos: 1.96201e+06 muA
** NormalTransistorNmos: 1.00031e+07 muA
** NormalTransistorPmos: -3.66389e+07 muA
** DiodeTransistorPmos: -1.48055e+08 muA
** DiodeTransistorPmos: -1.48055e+08 muA
** NormalTransistorNmos: 2.9611e+08 muA
** DiodeTransistorNmos: 2.96109e+08 muA
** NormalTransistorNmos: 1.48056e+08 muA
** NormalTransistorNmos: 1.48056e+08 muA
** NormalTransistorNmos: 1.70692e+08 muA
** NormalTransistorNmos: 1.70691e+08 muA
** NormalTransistorPmos: -1.70691e+08 muA
** NormalTransistorPmos: -1.7069e+08 muA
** NormalTransistorNmos: 1.7069e+08 muA
** NormalTransistorNmos: 1.70689e+08 muA
** NormalTransistorPmos: -1.70689e+08 muA
** NormalTransistorPmos: -1.7069e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 3.66381e+07 muA
** DiodeTransistorPmos: -1.96299e+06 muA
** DiodeTransistorPmos: -1.00039e+07 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.819001  V
** inOutputTransconductanceComplementarySecondStage: 3.78501  V
** inSourceTransconductanceComplementarySecondStage: 4.13301  V
** innerComplementarySecondStage: 0.567001  V
** inputVoltageBiasXXpXX0: 4.27001  V
** out: 2.5  V
** outFirstStage: 4.13301  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.34601  V
** innerStageBias: 0.168001  V
** innerTransconductance: 4.58901  V
** inner: 0.162001  V
** inner: 4.58901  V
** inner: 0.556001  V


.END