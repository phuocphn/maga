** Name: two_stage_single_output_op_amp_124_9

.MACRO two_stage_single_output_op_amp_124_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=8e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=128e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=99e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=393e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=7e-6
mTelescopicFirstStageLoad6 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=168e-6
mTelescopicFirstStageLoad7 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=168e-6
mMainBias8 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=165e-6
mTelescopicFirstStageLoad9 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=31e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=52e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=52e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=128e-6
mMainBias13 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=64e-6
mSecondStage1StageBias15 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=393e-6
mTelescopicFirstStageLoad16 outFirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=31e-6
mTelescopicFirstStageStageBias17 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=99e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=168e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=404e-6
mTelescopicFirstStageLoad20 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=5e-6 W=168e-6
mMainBias21 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=153e-6
mMainBias22 outVoltageBiasXXnXX3 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=37e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.2001e-12
.EOM two_stage_single_output_op_amp_124_9

** Expected Performance Values: 
** Gain: 146 dB
** Power consumption: 3.52301 mW
** Area: 11736 (mu_m)^2
** Transit frequency: 3.73201 MHz
** Transit frequency with error factor: 3.73202 MHz
** Slew rate: 5.08002 V/mu_s
** Phase margin: 60.1606°
** CMRR: 151 dB
** VoutMax: 4.63001 V
** VoutMin: 0.820001 V
** VcmMax: 3.76001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 7.88511e+07 muA
** NormalTransistorPmos: -7.42489e+07 muA
** NormalTransistorPmos: -1.76019e+07 muA
** NormalTransistorNmos: 1.98081e+07 muA
** NormalTransistorNmos: 1.98081e+07 muA
** DiodeTransistorPmos: -1.98089e+07 muA
** NormalTransistorPmos: -1.98099e+07 muA
** NormalTransistorPmos: -1.98089e+07 muA
** DiodeTransistorPmos: -1.98099e+07 muA
** NormalTransistorNmos: 5.72181e+07 muA
** DiodeTransistorNmos: 5.72171e+07 muA
** NormalTransistorNmos: 1.98091e+07 muA
** NormalTransistorNmos: 1.98091e+07 muA
** NormalTransistorNmos: 4.8419e+08 muA
** DiodeTransistorNmos: 4.84191e+08 muA
** NormalTransistorPmos: -4.84189e+08 muA
** DiodeTransistorNmos: 7.42481e+07 muA
** NormalTransistorNmos: 7.42471e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 1.76011e+07 muA
** DiodeTransistorPmos: -7.88519e+07 muA


** Expected Voltages: 
** ibias: 1.22801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.15201  V
** out: 2.5  V
** outFirstStage: 4.06801  V
** outInputVoltageBiasXXnXX1: 1.24601  V
** outSourceVoltageBiasXXnXX1: 0.623001  V
** outSourceVoltageBiasXXnXX2: 0.615001  V
** outVoltageBiasXXnXX3: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerOutputLoad2: 3.50801  V
** innerSourceLoad2: 4.25401  V
** innerTransistorStack1Load2: 4.25301  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.621001  V
** inner: 0.612001  V


.END