** Name: two_stage_single_output_op_amp_40_7

.MACRO two_stage_single_output_op_amp_40_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=150e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=26e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=23e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=5e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=26e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=150e-6
mMainBias10 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=323e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=5e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=190e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=23e-6
mMainBias16 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=479e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_40_7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 4.58301 mW
** Area: 2616 (mu_m)^2
** Transit frequency: 3.63701 MHz
** Transit frequency with error factor: 3.63206 MHz
** Slew rate: 8.34421 V/mu_s
** Phase margin: 63.5984°
** CMRR: 96 dB
** negPSRR: 92 dB
** posPSRR: 86 dB
** VoutMax: 4.25 V
** VoutMin: 0.220001 V
** VcmMax: 3.76001 V
** VcmMin: 1.54001 V


** Expected Currents: 
** NormalTransistorNmos: 1.20791e+07 muA
** NormalTransistorPmos: -2.13891e+08 muA
** DiodeTransistorPmos: -1.88089e+07 muA
** NormalTransistorPmos: -1.88079e+07 muA
** NormalTransistorPmos: -1.88069e+07 muA
** DiodeTransistorPmos: -1.88079e+07 muA
** NormalTransistorNmos: 3.76151e+07 muA
** DiodeTransistorNmos: 3.76141e+07 muA
** NormalTransistorNmos: 1.88081e+07 muA
** NormalTransistorNmos: 1.88081e+07 muA
** NormalTransistorNmos: 6.43049e+08 muA
** NormalTransistorPmos: -6.43048e+08 muA
** DiodeTransistorNmos: 2.13892e+08 muA
** NormalTransistorNmos: 2.13891e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.20799e+07 muA


** Expected Voltages: 
** ibias: 0.622001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.27801  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.17801  V
** outSourceVoltageBiasXXnXX1: 0.589001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.22301  V
** innerTransistorStack1Load1: 4.22401  V
** out1: 3.35801  V
** sourceTransconductance: 1.72901  V
** inner: 0.589001  V


.END