** Name: two_stage_single_output_op_amp_71_2

.MACRO two_stage_single_output_op_amp_71_2 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=53e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=18e-6
mSecondStage1StageBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=35e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=51e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=111e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=32e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=522e-6
mMainBias11 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=320e-6
mSecondStage1Transconductor12 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=148e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=53e-6
mMainBias14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=64e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerLoad2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=272e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=126e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=126e-6
mMainBias18 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=453e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=480e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=272e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.4001e-12
.EOM two_stage_single_output_op_amp_71_2

** Expected Performance Values: 
** Gain: 103 dB
** Power consumption: 5.17401 mW
** Area: 8499 (mu_m)^2
** Transit frequency: 4.47101 MHz
** Transit frequency with error factor: 4.46778 MHz
** Slew rate: 3.81869 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** VoutMax: 4.80001 V
** VoutMin: 0.310001 V
** VcmMax: 5.21001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 1.77684e+08 muA
** NormalTransistorNmos: 3.53631e+07 muA
** NormalTransistorPmos: -3.08003e+08 muA
** NormalTransistorPmos: -5.52339e+07 muA
** NormalTransistorPmos: -8.57099e+07 muA
** NormalTransistorPmos: -5.52339e+07 muA
** NormalTransistorPmos: -8.57099e+07 muA
** DiodeTransistorNmos: 5.52331e+07 muA
** NormalTransistorNmos: 5.52331e+07 muA
** NormalTransistorNmos: 6.09491e+07 muA
** NormalTransistorNmos: 6.09481e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 3.32422e+08 muA
** NormalTransistorNmos: 3.32421e+08 muA
** NormalTransistorPmos: -3.32421e+08 muA
** DiodeTransistorNmos: 3.08004e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.77683e+08 muA
** DiodeTransistorPmos: -3.53639e+07 muA


** Expected Voltages: 
** ibias: 0.633001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.983001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXpXX2: 4.24001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.562001  V
** innerStageBias: 0.428001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 0.415001  V


.END