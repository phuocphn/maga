** Name: two_stage_single_output_op_amp_9_8

.MACRO two_stage_single_output_op_amp_9_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=51e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=9e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=9e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=23e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=344e-6
mSecondStage1StageBias8 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=333e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=9e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mSimpleFirstStageLoad11 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=51e-6
mMainBias12 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=18e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=56e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=8e-6 W=124e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_9_8

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 3.22801 mW
** Area: 4357 (mu_m)^2
** Transit frequency: 2.97301 MHz
** Transit frequency with error factor: 2.96853 MHz
** Slew rate: 8.32151 V/mu_s
** Phase margin: 65.3172°
** CMRR: 95 dB
** negPSRR: 93 dB
** posPSRR: 85 dB
** VoutMax: 4.25 V
** VoutMin: 0.480001 V
** VcmMax: 4.17001 V
** VcmMin: 1.05001 V


** Expected Currents: 
** NormalTransistorNmos: 9.88301e+06 muA
** NormalTransistorPmos: -1.93919e+07 muA
** NormalTransistorPmos: -1.88939e+07 muA
** NormalTransistorPmos: -1.88939e+07 muA
** DiodeTransistorPmos: -1.88939e+07 muA
** NormalTransistorNmos: 3.77871e+07 muA
** NormalTransistorNmos: 1.88931e+07 muA
** NormalTransistorNmos: 1.88931e+07 muA
** NormalTransistorNmos: 5.6859e+08 muA
** NormalTransistorNmos: 5.68589e+08 muA
** NormalTransistorPmos: -5.68589e+08 muA
** DiodeTransistorNmos: 1.93911e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.88399e+06 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.886001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 3.69601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.02901  V
** out1: 3.20501  V
** sourceTransconductance: 1.64801  V
** innerStageBias: 0.198001  V


.END