** Name: two_stage_single_output_op_amp_80_10

.MACRO two_stage_single_output_op_amp_80_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=26e-6
mMainBias2 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=9e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=56e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mMainBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=10e-6 W=459e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=55e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=55e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=31e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=31e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=56e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias14 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mSecondStage1StageBias15 out inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=397e-6
mFoldedCascodeFirstStageLoad16 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=459e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=137e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=370e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=370e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=547e-6
mMainBias21 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=130e-6
mMainBias22 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=67e-6
mSecondStage1Transconductor23 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad24 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=137e-6
mMainBias25 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.4001e-12
.EOM two_stage_single_output_op_amp_80_10

** Expected Performance Values: 
** Gain: 132 dB
** Power consumption: 10.2811 mW
** Area: 14812 (mu_m)^2
** Transit frequency: 8.625 MHz
** Transit frequency with error factor: 8.62522 MHz
** Slew rate: 8.12912 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.510001 V
** VcmMax: 5.24001 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorNmos: 1.11687e+08 muA
** NormalTransistorPmos: -2.52449e+07 muA
** NormalTransistorPmos: -6.19079e+07 muA
** NormalTransistorPmos: -3.23169e+07 muA
** NormalTransistorPmos: -1.18088e+08 muA
** NormalTransistorPmos: -1.77131e+08 muA
** NormalTransistorPmos: -1.18092e+08 muA
** NormalTransistorPmos: -1.77137e+08 muA
** NormalTransistorNmos: 1.18091e+08 muA
** NormalTransistorNmos: 1.18092e+08 muA
** NormalTransistorNmos: 1.18093e+08 muA
** NormalTransistorNmos: 1.18092e+08 muA
** NormalTransistorNmos: 1.18088e+08 muA
** DiodeTransistorNmos: 1.18087e+08 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorNmos: 1.45079e+09 muA
** NormalTransistorPmos: -1.45078e+09 muA
** NormalTransistorPmos: -1.45078e+09 muA
** DiodeTransistorNmos: 2.52441e+07 muA
** NormalTransistorNmos: 2.52431e+07 muA
** DiodeTransistorNmos: 6.19071e+07 muA
** DiodeTransistorNmos: 3.23161e+07 muA
** DiodeTransistorPmos: -1.11686e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.938001  V
** inputVoltageBiasXXnXX3: 0.912001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.05201  V
** outInputVoltageBiasXXnXX1: 1.12601  V
** outSourceVoltageBiasXXnXX1: 0.563001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.564001  V
** innerTransistorStack1Load2: 0.358001  V
** innerTransistorStack2Load2: 0.359001  V
** sourceGCC1: 4.46901  V
** sourceGCC2: 4.46901  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.61601  V
** inner: 0.563001  V


.END