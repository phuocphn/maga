** Name: two_stage_single_output_op_amp_86_1

.MACRO two_stage_single_output_op_amp_86_1 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=84e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=524e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=8e-6 W=58e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=84e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=264e-6
mTelescopicFirstStageLoad7 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=14e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=555e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=8e-6 W=8e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=142e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=142e-6
mSecondStage1StageBias12 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=238e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=8e-6 W=8e-6
mMainBias14 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=185e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=230e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.90001e-12
.EOM two_stage_single_output_op_amp_86_1

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 5.60601 mW
** Area: 10556 (mu_m)^2
** Transit frequency: 3.15901 MHz
** Transit frequency with error factor: 3.1586 MHz
** Slew rate: 13.2743 V/mu_s
** Phase margin: 60.1606°
** CMRR: 118 dB
** VoutMax: 4.57001 V
** VoutMin: 0.300001 V
** VcmMax: 3.73001 V
** VcmMin: 1.37001 V


** Expected Currents: 
** NormalTransistorNmos: 3.35017e+08 muA
** NormalTransistorPmos: -3.14491e+08 muA
** NormalTransistorPmos: -2.66659e+07 muA
** NormalTransistorPmos: -2.66659e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** DiodeTransistorNmos: 2.66651e+07 muA
** NormalTransistorPmos: -3.88351e+08 muA
** NormalTransistorPmos: -2.66669e+07 muA
** NormalTransistorPmos: -2.66669e+07 muA
** NormalTransistorNmos: 3.98276e+08 muA
** NormalTransistorPmos: -3.98275e+08 muA
** DiodeTransistorNmos: 3.14492e+08 muA
** DiodeTransistorPmos: -3.35016e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.00201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outVoltageBiasXXnXX0: 0.574001  V
** outVoltageBiasXXpXX1: 1.17001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.33401  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 2.96101  V
** sourceGCC2: 2.96101  V


.END