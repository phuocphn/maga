** Name: two_stage_single_output_op_amp_113_12

.MACRO two_stage_single_output_op_amp_113_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=2e-6 W=6e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=82e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=394e-6
mMainBias4 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=198e-6
mTelescopicFirstStageLoad6 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=73e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad9 FirstStageYinnerLoad2 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=40e-6
mTelescopicFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=558e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=121e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=121e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=82e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mSecondStage1StageBias15 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=394e-6
mTelescopicFirstStageLoad16 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=40e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=35e-6
mTelescopicFirstStageStageBias18 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=168e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=390e-6
mMainBias20 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=13e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mTelescopicFirstStageLoad22 outFirstStage FirstStageYinnerLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=73e-6
mMainBias23 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=118e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20e-12
.EOM two_stage_single_output_op_amp_113_12

** Expected Performance Values: 
** Gain: 150 dB
** Power consumption: 4.69401 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 2.71301 MHz
** Transit frequency with error factor: 2.71154 MHz
** Slew rate: 6.75812 V/mu_s
** Phase margin: 60.1606°
** CMRR: 85 dB
** VoutMax: 4.64001 V
** VoutMin: 0.940001 V
** VcmMax: 4.49001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorNmos: 1.70131e+07 muA
** NormalTransistorNmos: 3.50271e+07 muA
** NormalTransistorPmos: -5.58819e+07 muA
** NormalTransistorPmos: -4.97843e+08 muA
** NormalTransistorNmos: 2.56061e+07 muA
** NormalTransistorNmos: 2.56061e+07 muA
** DiodeTransistorPmos: -2.56069e+07 muA
** NormalTransistorPmos: -2.56069e+07 muA
** NormalTransistorNmos: 5.49057e+08 muA
** NormalTransistorNmos: 5.49056e+08 muA
** NormalTransistorNmos: 2.56071e+07 muA
** NormalTransistorNmos: 2.56071e+07 muA
** NormalTransistorNmos: 2.71803e+08 muA
** DiodeTransistorNmos: 2.71802e+08 muA
** NormalTransistorPmos: -2.71802e+08 muA
** NormalTransistorPmos: -2.71803e+08 muA
** DiodeTransistorNmos: 5.58811e+07 muA
** NormalTransistorNmos: 5.58801e+07 muA
** DiodeTransistorNmos: 4.97844e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.70139e+07 muA
** DiodeTransistorPmos: -3.50279e+07 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.35001  V
** inputVoltageBiasXXpXX0: 3.46001  V
** out: 2.5  V
** outFirstStage: 4.23801  V
** outSourceVoltageBiasXXnXX1: 0.675001  V
** outSourceVoltageBiasXXnXX3: 0.558001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX1: 3.99201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerLoad2: 4.23701  V
** innerStageBias: 0.477001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.71501  V
** inner: 0.675001  V


.END