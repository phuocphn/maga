** Name: two_stage_single_output_op_amp_204_9

.MACRO two_stage_single_output_op_amp_204_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=6e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=83e-6
mMainBias4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=11e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=52e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=535e-6
mMainBias7 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=48e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=11e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=52e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=83e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=535e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=6e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=11e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=264e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=333e-6
mSimpleFirstStageLoad18 outFirstStage ibias sourcePmos sourcePmos pmos4 L=4e-6 W=264e-6
mMainBias19 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=315e-6
mMainBias20 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=161e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.60001e-12
.EOM two_stage_single_output_op_amp_204_9

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 9.61001 mW
** Area: 9396 (mu_m)^2
** Transit frequency: 6.66901 MHz
** Transit frequency with error factor: 6.6561 MHz
** Slew rate: 6.28502 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 1.07001 V
** VcmMax: 5.19001 V
** VcmMin: 1.35001 V


** Expected Currents: 
** NormalTransistorPmos: -6.61299e+07 muA
** NormalTransistorPmos: -3.42109e+07 muA
** DiodeTransistorNmos: 3.46511e+07 muA
** NormalTransistorNmos: 3.46521e+07 muA
** NormalTransistorNmos: 3.46511e+07 muA
** DiodeTransistorNmos: 3.46521e+07 muA
** NormalTransistorPmos: -5.56029e+07 muA
** NormalTransistorPmos: -5.56029e+07 muA
** NormalTransistorNmos: 4.19011e+07 muA
** DiodeTransistorNmos: 4.19001e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 1.69055e+09 muA
** DiodeTransistorNmos: 1.69055e+09 muA
** NormalTransistorPmos: -1.69054e+09 muA
** DiodeTransistorNmos: 6.61291e+07 muA
** NormalTransistorNmos: 6.61301e+07 muA
** DiodeTransistorNmos: 3.42101e+07 muA
** NormalTransistorNmos: 3.42091e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.20001  V
** outInputVoltageBiasXXnXX2: 1.47601  V
** outSourceVoltageBiasXXnXX1: 0.600001  V
** outSourceVoltageBiasXXnXX2: 0.738001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.04801  V
** innerTransistorStack1Load1: 1.04801  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 0.601001  V
** inner: 0.738001  V


.END