** Name: two_stage_single_output_op_amp_48_5

.MACRO two_stage_single_output_op_amp_48_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=6e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=95e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=10e-6 W=95e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=35e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=486e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=180e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=13e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=41e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=41e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=176e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=13e-6
mMainBias13 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=54e-6
mMainBias14 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=82e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=95e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=99e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=99e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=62e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=35e-6
mSecondStage1StageBias20 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=486e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=10e-6 W=95e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_48_5

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 4.85401 mW
** Area: 8048 (mu_m)^2
** Transit frequency: 4.88601 MHz
** Transit frequency with error factor: 4.88544 MHz
** Slew rate: 5.88417 V/mu_s
** Phase margin: 66.4632°
** CMRR: 133 dB
** VoutMax: 3.85001 V
** VoutMin: 0.550001 V
** VcmMax: 3.89001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 5.35251e+07 muA
** NormalTransistorNmos: 8.04411e+07 muA
** NormalTransistorNmos: 2.66081e+07 muA
** NormalTransistorNmos: 4.02211e+07 muA
** NormalTransistorNmos: 2.66081e+07 muA
** NormalTransistorNmos: 4.02211e+07 muA
** DiodeTransistorPmos: -2.66089e+07 muA
** NormalTransistorPmos: -2.66099e+07 muA
** NormalTransistorPmos: -2.66089e+07 muA
** DiodeTransistorPmos: -2.66099e+07 muA
** NormalTransistorPmos: -2.72289e+07 muA
** NormalTransistorPmos: -1.36139e+07 muA
** NormalTransistorPmos: -1.36139e+07 muA
** NormalTransistorNmos: 7.46399e+08 muA
** NormalTransistorPmos: -7.46398e+08 muA
** DiodeTransistorPmos: -7.46399e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.35259e+07 muA
** NormalTransistorPmos: -5.35269e+07 muA
** DiodeTransistorPmos: -8.04419e+07 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.956001  V
** outInputVoltageBiasXXpXX1: 3.28401  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.14201  V
** outVoltageBiasXXpXX2: 4.08401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.10401  V
** innerTransistorStack1Load2: 4.10101  V
** out1: 3.14301  V
** sourceGCC1: 0.535001  V
** sourceGCC2: 0.535001  V
** sourceTransconductance: 3.26001  V
** inner: 4.14001  V


.END