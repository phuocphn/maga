** Name: two_stage_single_output_op_amp_65_10

.MACRO two_stage_single_output_op_amp_65_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=124e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=59e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=38e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=38e-6
mSecondStage1StageBias8 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=336e-6
mFoldedCascodeFirstStageLoad9 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=59e-6
mMainBias10 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=63e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=600e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=102e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=22e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=22e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=57e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=581e-6
mMainBias19 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=262e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=558e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=102e-6
mMainBias22 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=570e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.90001e-12
.EOM two_stage_single_output_op_amp_65_10

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 4.98901 mW
** Area: 14997 (mu_m)^2
** Transit frequency: 5.25901 MHz
** Transit frequency with error factor: 5.25905 MHz
** Slew rate: 8.25087 V/mu_s
** Phase margin: 60.1606°
** CMRR: 136 dB
** VoutMax: 4.25 V
** VoutMin: 0.150001 V
** VcmMax: 3.23001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorPmos: -4.56759e+07 muA
** NormalTransistorPmos: -2.10219e+07 muA
** NormalTransistorNmos: 4.90231e+07 muA
** NormalTransistorNmos: 7.35331e+07 muA
** NormalTransistorNmos: 4.90251e+07 muA
** NormalTransistorNmos: 7.35351e+07 muA
** NormalTransistorPmos: -4.90239e+07 muA
** NormalTransistorPmos: -4.90249e+07 muA
** NormalTransistorPmos: -4.90259e+07 muA
** NormalTransistorPmos: -4.90249e+07 muA
** NormalTransistorPmos: -4.90219e+07 muA
** NormalTransistorPmos: -4.90209e+07 muA
** NormalTransistorPmos: -2.45109e+07 muA
** NormalTransistorPmos: -2.45109e+07 muA
** NormalTransistorNmos: 6.42096e+08 muA
** NormalTransistorPmos: -6.42095e+08 muA
** NormalTransistorPmos: -6.42096e+08 muA
** DiodeTransistorNmos: 4.56751e+07 muA
** DiodeTransistorNmos: 2.10211e+07 muA
** DiodeTransistorPmos: -1.21839e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.556001  V
** out: 2.5  V
** outFirstStage: 3.93901  V
** outVoltageBiasXXnXX1: 0.927001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.46901  V
** innerTransistorStack1Load2: 4.41401  V
** innerTransistorStack2Load2: 4.41401  V
** out1: 4.09701  V
** sourceGCC1: 0.351001  V
** sourceGCC2: 0.351001  V
** sourceTransconductance: 3.31301  V
** innerTransconductance: 4.50301  V


.END