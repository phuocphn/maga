** Name: two_stage_single_output_op_amp_190_9

.MACRO two_stage_single_output_op_amp_190_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=7e-6 W=10e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=155e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=1e-6 W=12e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=86e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=368e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=13e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=74e-6
mSimpleFirstStageLoad9 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=7e-6 W=10e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=86e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=155e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=368e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=20e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=74e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=51e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=51e-6
mSimpleFirstStageLoad18 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=66e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=111e-6
mSimpleFirstStageLoad20 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=66e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=37e-6
mMainBias22 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=22e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.60001e-12
.EOM two_stage_single_output_op_amp_190_9

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 7.09601 mW
** Area: 5369 (mu_m)^2
** Transit frequency: 4.32601 MHz
** Transit frequency with error factor: 4.32337 MHz
** Slew rate: 4.07662 V/mu_s
** Phase margin: 60.1606°
** CMRR: 110 dB
** VoutMax: 4.25 V
** VoutMin: 0.780001 V
** VcmMax: 4.59001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorPmos: -6.28979e+07 muA
** NormalTransistorPmos: -3.70419e+07 muA
** NormalTransistorNmos: 6.85401e+07 muA
** NormalTransistorNmos: 6.85411e+07 muA
** DiodeTransistorNmos: 6.85401e+07 muA
** NormalTransistorPmos: -8.61589e+07 muA
** NormalTransistorPmos: -8.61599e+07 muA
** NormalTransistorPmos: -8.61599e+07 muA
** NormalTransistorPmos: -8.61599e+07 muA
** NormalTransistorNmos: 3.52351e+07 muA
** DiodeTransistorNmos: 3.52341e+07 muA
** NormalTransistorNmos: 1.76181e+07 muA
** NormalTransistorNmos: 1.76181e+07 muA
** NormalTransistorNmos: 1.12703e+09 muA
** DiodeTransistorNmos: 1.12703e+09 muA
** NormalTransistorPmos: -1.12702e+09 muA
** DiodeTransistorNmos: 6.28971e+07 muA
** NormalTransistorNmos: 6.28961e+07 muA
** DiodeTransistorNmos: 3.70411e+07 muA
** NormalTransistorNmos: 3.70401e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.14401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.12001  V
** outInputVoltageBiasXXnXX2: 1.19001  V
** outSourceVoltageBiasXXnXX1: 0.560001  V
** outSourceVoltageBiasXXnXX2: 0.595001  V
** outSourceVoltageBiasXXpXX1: 4.00201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.08901  V
** innerTransistorStack2Load1: 1.15501  V
** innerTransistorStack2Load2: 4.08901  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 0.560001  V
** inner: 0.594001  V


.END