** Name: two_stage_single_output_op_amp_188_10

.MACRO two_stage_single_output_op_amp_188_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=63e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=25e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=27e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=61e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=69e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=28e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=63e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=61e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=27e-6
mMainBias11 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=271e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=9e-6 W=600e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=1e-6 W=14e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=28e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=306e-6
mSimpleFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=230e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=394e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=523e-6
mSimpleFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=230e-6
mMainBias20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.20001e-12
.EOM two_stage_single_output_op_amp_188_10

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 5.99701 mW
** Area: 14834 (mu_m)^2
** Transit frequency: 4.56001 MHz
** Transit frequency with error factor: 4.49614 MHz
** Slew rate: 4.29797 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.66001 V
** VoutMin: 0.210001 V
** VcmMax: 5.11001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorNmos: 1.07654e+08 muA
** NormalTransistorPmos: -1.56019e+07 muA
** NormalTransistorNmos: 3.35847e+08 muA
** NormalTransistorNmos: 3.35848e+08 muA
** DiodeTransistorNmos: 3.35847e+08 muA
** NormalTransistorPmos: -3.53623e+08 muA
** NormalTransistorPmos: -3.53623e+08 muA
** NormalTransistorNmos: 3.55531e+07 muA
** DiodeTransistorNmos: 3.55521e+07 muA
** NormalTransistorNmos: 1.77771e+07 muA
** NormalTransistorNmos: 1.77771e+07 muA
** NormalTransistorNmos: 2.37111e+08 muA
** NormalTransistorPmos: -2.3711e+08 muA
** NormalTransistorPmos: -2.37111e+08 muA
** DiodeTransistorNmos: 1.56011e+07 muA
** NormalTransistorNmos: 1.56001e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.21839e+08 muA
** DiodeTransistorPmos: -1.07653e+08 muA


** Expected Voltages: 
** ibias: 0.611001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.14201  V
** out: 2.5  V
** outFirstStage: 4.25201  V
** outInputVoltageBiasXXnXX1: 1.24801  V
** outSourceVoltageBiasXXnXX1: 0.624001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.40901  V
** inner: 0.624001  V


.END