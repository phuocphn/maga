** Name: two_stage_single_output_op_amp_54_6

.MACRO two_stage_single_output_op_amp_54_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=35e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=8e-6 W=38e-6
mMainBias4 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=5e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=541e-6
mMainBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=31e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=20e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=70e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=70e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=34e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=34e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=94e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=74e-6
mSecondStage1Transconductor14 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=570e-6
mFoldedCascodeFirstStageLoad15 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=20e-6
mMainBias16 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=138e-6
mMainBias17 outInputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=83e-6
mFoldedCascodeFirstStageLoad18 FirstStageYinnerSourceLoad2 outInputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=61e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=43e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=43e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=38e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=8e-6 W=541e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outInputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=61e-6
mMainBias24 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=83e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_54_6

** Expected Performance Values: 
** Gain: 174 dB
** Power consumption: 3.71501 mW
** Area: 14994 (mu_m)^2
** Transit frequency: 6.13301 MHz
** Transit frequency with error factor: 6.13312 MHz
** Slew rate: 4.21477 V/mu_s
** Phase margin: 62.4525°
** CMRR: 146 dB
** VoutMax: 3.09001 V
** VoutMin: 0.440001 V
** VcmMax: 5.11001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorNmos: 3.86791e+07 muA
** NormalTransistorNmos: 2.36901e+07 muA
** NormalTransistorPmos: -6.34339e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -3.22219e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -3.22219e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 2.63471e+07 muA
** NormalTransistorNmos: 1.31731e+07 muA
** NormalTransistorNmos: 1.31731e+07 muA
** NormalTransistorNmos: 5.4282e+08 muA
** NormalTransistorNmos: 5.42819e+08 muA
** NormalTransistorPmos: -5.42819e+08 muA
** DiodeTransistorPmos: -5.4282e+08 muA
** DiodeTransistorNmos: 6.34331e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.86799e+07 muA
** NormalTransistorPmos: -3.86809e+07 muA
** DiodeTransistorPmos: -2.36909e+07 muA
** DiodeTransistorPmos: -2.36919e+07 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.700001  V
** outInputVoltageBiasXXpXX1: 2.52601  V
** outInputVoltageBiasXXpXX2: 2.85001  V
** outSourceVoltageBiasXXpXX1: 3.76301  V
** outSourceVoltageBiasXXpXX2: 4.14501  V
** outVoltageBiasXXnXX1: 0.905001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.350001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 3.60101  V
** sourceGCC2: 3.60101  V
** sourceTransconductance: 1.94301  V
** innerTransconductance: 0.350001  V
** inner: 3.76201  V


.END