** Name: two_stage_single_output_op_amp_38_7

.MACRO two_stage_single_output_op_amp_38_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=16e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=56e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=132e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=34e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=56e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=16e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=34e-6
mMainBias11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=135e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=61e-6
mSimpleFirstStageLoad13 FirstStageYinnerSourceLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=107e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=22e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=22e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=579e-6
mSimpleFirstStageLoad17 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=107e-6
mMainBias18 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=12e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_38_7

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 4.30401 mW
** Area: 6241 (mu_m)^2
** Transit frequency: 4.95701 MHz
** Transit frequency with error factor: 4.95407 MHz
** Slew rate: 4.67171 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 105 dB
** posPSRR: 99 dB
** VoutMax: 4.58001 V
** VoutMin: 0.150001 V
** VcmMax: 4.88001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 1.34024e+08 muA
** NormalTransistorNmos: 6.09191e+07 muA
** NormalTransistorPmos: -1.21839e+07 muA
** NormalTransistorPmos: -2.15869e+07 muA
** NormalTransistorPmos: -2.15879e+07 muA
** NormalTransistorPmos: -2.15869e+07 muA
** NormalTransistorPmos: -2.15879e+07 muA
** NormalTransistorNmos: 4.31711e+07 muA
** DiodeTransistorNmos: 4.31701e+07 muA
** NormalTransistorNmos: 2.15861e+07 muA
** NormalTransistorNmos: 2.15861e+07 muA
** NormalTransistorNmos: 6.00477e+08 muA
** NormalTransistorPmos: -6.00476e+08 muA
** DiodeTransistorNmos: 1.21831e+07 muA
** NormalTransistorNmos: 1.21821e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.34023e+08 muA
** DiodeTransistorPmos: -6.09199e+07 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.01701  V
** outInputVoltageBiasXXnXX1: 1.19001  V
** outSourceVoltageBiasXXnXX1: 0.595001  V
** outVoltageBiasXXpXX0: 3.68601  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.91201  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94501  V
** inner: 0.595001  V


.END