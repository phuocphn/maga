** Name: two_stage_single_output_op_amp_152_9

.MACRO two_stage_single_output_op_amp_152_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=8e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=7e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=272e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=10e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=58e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=272e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=8e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=58e-6
mSimpleFirstStageLoad15 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=26e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=35e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=35e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=175e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=26e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=32e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_152_9

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 9.82901 mW
** Area: 5879 (mu_m)^2
** Transit frequency: 5.18201 MHz
** Transit frequency with error factor: 5.17997 MHz
** Slew rate: 4.88341 V/mu_s
** Phase margin: 68.182°
** CMRR: 108 dB
** VoutMax: 4.25 V
** VoutMin: 1.87001 V
** VcmMax: 4.54001 V
** VcmMin: 0.890001 V


** Expected Currents: 
** NormalTransistorPmos: -4.58169e+07 muA
** NormalTransistorPmos: -2.17689e+07 muA
** DiodeTransistorNmos: 3.96021e+07 muA
** NormalTransistorNmos: 3.96031e+07 muA
** NormalTransistorNmos: 3.96021e+07 muA
** DiodeTransistorNmos: 3.96031e+07 muA
** NormalTransistorPmos: -5.06499e+07 muA
** NormalTransistorPmos: -5.06509e+07 muA
** NormalTransistorPmos: -5.06499e+07 muA
** NormalTransistorPmos: -5.06509e+07 muA
** NormalTransistorNmos: 2.20931e+07 muA
** NormalTransistorNmos: 1.10471e+07 muA
** NormalTransistorNmos: 1.10471e+07 muA
** NormalTransistorNmos: 1.77685e+09 muA
** DiodeTransistorNmos: 1.77685e+09 muA
** NormalTransistorPmos: -1.77684e+09 muA
** DiodeTransistorNmos: 4.58161e+07 muA
** NormalTransistorNmos: 4.58151e+07 muA
** DiodeTransistorNmos: 2.17681e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 2.27401  V
** outSourceVoltageBiasXXnXX1: 1.13701  V
** outSourceVoltageBiasXXpXX1: 4.03501  V
** outVoltageBiasXXnXX2: 0.738001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerTransistorStack1Load1: 1.04801  V
** innerTransistorStack1Load2: 4.16401  V
** innerTransistorStack2Load1: 1.04801  V
** innerTransistorStack2Load2: 4.16401  V
** sourceTransconductance: 1.94501  V
** inner: 1.13001  V


.END