** Name: two_stage_single_output_op_amp_54_1

.MACRO two_stage_single_output_op_amp_54_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=10e-6 W=37e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=16e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=46e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=121e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=65e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=65e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=15e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=15e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=10e-6 W=214e-6
mMainBias11 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=490e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=121e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=121e-6
mMainBias14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=235e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=106e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=53e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=53e-6
mMainBias18 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=36e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=580e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=106e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.70001e-12
.EOM two_stage_single_output_op_amp_54_1

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 5.97001 mW
** Area: 14635 (mu_m)^2
** Transit frequency: 6.20801 MHz
** Transit frequency with error factor: 6.20823 MHz
** Slew rate: 4.40839 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.61001 V
** VoutMin: 0.390001 V
** VcmMax: 5.02001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorNmos: 1.31994e+08 muA
** NormalTransistorNmos: 6.31451e+07 muA
** NormalTransistorPmos: -4.94179e+07 muA
** NormalTransistorPmos: -4.30499e+07 muA
** NormalTransistorPmos: -7.16209e+07 muA
** NormalTransistorPmos: -4.30499e+07 muA
** NormalTransistorPmos: -7.16209e+07 muA
** NormalTransistorNmos: 4.30491e+07 muA
** NormalTransistorNmos: 4.30481e+07 muA
** NormalTransistorNmos: 4.30491e+07 muA
** NormalTransistorNmos: 4.30481e+07 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 7.96189e+08 muA
** NormalTransistorPmos: -7.96188e+08 muA
** DiodeTransistorNmos: 4.94171e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.31993e+08 muA
** DiodeTransistorPmos: -6.31459e+07 muA


** Expected Voltages: 
** ibias: 0.583001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.976001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.798001  V
** outVoltageBiasXXpXX2: 4.04601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.582001  V
** innerTransistorStack1Load2: 0.376001  V
** innerTransistorStack2Load2: 0.377001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V


.END