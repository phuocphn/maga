** Name: symmetrical_op_amp150

.MACRO symmetrical_op_amp150 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias2 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=189e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=101e-6
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=101e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=93e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=93e-6
mSymmetricalFirstStageLoad10 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=153e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=4e-6 W=115e-6
mSecondStage1Transconductor12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=115e-6
mSymmetricalFirstStageLoad13 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=153e-6
mSymmetricalFirstStageStageBias14 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=189e-6
mSecondStage1StageBias15 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mSymmetricalFirstStageTransconductor17 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=567e-6
mSecondStage1StageBias18 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=185e-6
mSymmetricalFirstStageTransconductor19 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=567e-6
mMainBias20 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp150

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 2.01001 mW
** Area: 8583 (mu_m)^2
** Transit frequency: 7.21101 MHz
** Transit frequency with error factor: 7.21147 MHz
** Slew rate: 8.82469 V/mu_s
** Phase margin: 80.2142°
** CMRR: 152 dB
** negPSRR: 51 dB
** posPSRR: 69 dB
** VoutMax: 3.94001 V
** VoutMin: 0.340001 V
** VcmMax: 3 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.22259e+07 muA
** NormalTransistorNmos: 9.62871e+07 muA
** NormalTransistorNmos: 9.62861e+07 muA
** NormalTransistorNmos: 9.62871e+07 muA
** NormalTransistorNmos: 9.62861e+07 muA
** NormalTransistorPmos: -1.92574e+08 muA
** DiodeTransistorPmos: -1.92573e+08 muA
** NormalTransistorPmos: -9.62879e+07 muA
** NormalTransistorPmos: -9.62879e+07 muA
** NormalTransistorNmos: 8.85651e+07 muA
** NormalTransistorNmos: 8.85661e+07 muA
** NormalTransistorPmos: -8.85659e+07 muA
** NormalTransistorPmos: -8.85669e+07 muA
** DiodeTransistorPmos: -8.85679e+07 muA
** DiodeTransistorPmos: -8.85689e+07 muA
** NormalTransistorNmos: 8.85671e+07 muA
** NormalTransistorNmos: 8.85661e+07 muA
** DiodeTransistorNmos: 1.22251e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.19701  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 4.10701  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 2.83601  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.745001  V
** outSourceVoltageBiasXXpXX1: 4.10001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.167001  V
** innerTransistorStack2Load1: 0.167001  V
** sourceTransconductance: 3.25801  V
** innerStageBias: 3.56301  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V
** inner: 4.09401  V


.END