** Name: two_stage_single_output_op_amp_187_10

.MACRO two_stage_single_output_op_amp_187_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=199e-6
mSecondStage1StageBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=504e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=42e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=110e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=60e-6
mSecondStage1StageBias10 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=546e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=16e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=110e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=486e-6
mMainBias14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=517e-6
mSimpleFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=218e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=519e-6
mMainBias17 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=537e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=480e-6
mSimpleFirstStageLoad19 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=218e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.5e-12
.EOM two_stage_single_output_op_amp_187_10

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 12.5341 mW
** Area: 13894 (mu_m)^2
** Transit frequency: 5.86101 MHz
** Transit frequency with error factor: 5.81484 MHz
** Slew rate: 5.52351 V/mu_s
** Phase margin: 60.1606°
** CMRR: 95 dB
** VoutMax: 4.41001 V
** VoutMin: 0.150001 V
** VcmMax: 4.93001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 4.7721e+08 muA
** NormalTransistorNmos: 5.08841e+08 muA
** NormalTransistorPmos: -5.42157e+08 muA
** NormalTransistorNmos: 1.95517e+08 muA
** NormalTransistorNmos: 1.95518e+08 muA
** DiodeTransistorNmos: 1.95517e+08 muA
** NormalTransistorPmos: -2.16467e+08 muA
** NormalTransistorPmos: -2.16467e+08 muA
** NormalTransistorNmos: 4.19011e+07 muA
** NormalTransistorNmos: 4.19001e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 5.35614e+08 muA
** NormalTransistorPmos: -5.35613e+08 muA
** NormalTransistorPmos: -5.35614e+08 muA
** DiodeTransistorNmos: 5.42158e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.77209e+08 muA
** DiodeTransistorPmos: -5.0884e+08 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.715001  V
** out: 2.5  V
** outFirstStage: 4.09501  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 3.96301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.153001  V
** innerTransistorStack2Load1: 1.15001  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.49901  V


.END