** Name: two_stage_single_output_op_amp_147_12

.MACRO two_stage_single_output_op_amp_147_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=5e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=10e-6 W=34e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=6e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=322e-6
mSecondStage1StageBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=90e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=10e-6 W=389e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mMainBias12 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=447e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=322e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=5e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=90e-6
mMainBias16 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=26e-6
mSimpleFirstStageLoad17 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=57e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=483e-6
mSecondStage1Transconductor19 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad20 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=57e-6
mMainBias21 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=13e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.4001e-12
.EOM two_stage_single_output_op_amp_147_12

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 8.75301 mW
** Area: 14979 (mu_m)^2
** Transit frequency: 6.95401 MHz
** Transit frequency with error factor: 6.94384 MHz
** Slew rate: 6.55376 V/mu_s
** Phase margin: 60.1606°
** CMRR: 86 dB
** VoutMax: 4.25 V
** VoutMin: 1.49001 V
** VcmMax: 4.84001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorNmos: 1.31994e+08 muA
** NormalTransistorNmos: 7.54801e+06 muA
** NormalTransistorPmos: -2.49689e+07 muA
** DiodeTransistorNmos: 5.22821e+07 muA
** DiodeTransistorNmos: 5.22831e+07 muA
** NormalTransistorNmos: 5.22821e+07 muA
** NormalTransistorNmos: 5.22831e+07 muA
** NormalTransistorPmos: -1.09421e+08 muA
** NormalTransistorPmos: -1.09421e+08 muA
** NormalTransistorNmos: 1.14278e+08 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 1.35721e+09 muA
** DiodeTransistorNmos: 1.35721e+09 muA
** NormalTransistorPmos: -1.3572e+09 muA
** NormalTransistorPmos: -1.35721e+09 muA
** DiodeTransistorNmos: 2.49681e+07 muA
** NormalTransistorNmos: 2.49671e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.31993e+08 muA
** DiodeTransistorPmos: -7.54899e+06 muA


** Expected Voltages: 
** ibias: 0.591001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.04001  V
** outInputVoltageBiasXXnXX1: 1.89801  V
** outSourceVoltageBiasXXnXX1: 0.949001  V
** outVoltageBiasXXpXX2: 3.87101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.10501  V
** innerSourceLoad1: 1.08901  V
** innerTransistorStack2Load1: 1.08901  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.60401  V
** inner: 0.948001  V


.END