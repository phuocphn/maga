** Name: two_stage_single_output_op_amp_76_8

.MACRO two_stage_single_output_op_amp_76_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=56e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=463e-6
mFoldedCascodeFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=167e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=50e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=110e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=56e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=5e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=5e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=167e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=380e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=463e-6
mSecondStage1StageBias14 out outVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=390e-6
mFoldedCascodeFirstStageLoad15 outFirstStage outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=20e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=54e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=91e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=91e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=261e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=54e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=208e-6
mMainBias22 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=597e-6
mMainBias23 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=251e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_76_8

** Expected Performance Values: 
** Gain: 112 dB
** Power consumption: 10.7901 mW
** Area: 13114 (mu_m)^2
** Transit frequency: 4.01701 MHz
** Transit frequency with error factor: 4.01683 MHz
** Slew rate: 11.9099 V/mu_s
** Phase margin: 67.6091°
** CMRR: 130 dB
** VoutMax: 4.25 V
** VoutMin: 0.450001 V
** VcmMax: 5.17001 V
** VcmMin: 1.88001 V


** Expected Currents: 
** NormalTransistorPmos: -2.10885e+08 muA
** NormalTransistorPmos: -6.04793e+08 muA
** NormalTransistorPmos: -2.54482e+08 muA
** NormalTransistorPmos: -5.38289e+07 muA
** NormalTransistorPmos: -9.22619e+07 muA
** NormalTransistorPmos: -5.38289e+07 muA
** NormalTransistorPmos: -9.22619e+07 muA
** DiodeTransistorNmos: 5.38281e+07 muA
** NormalTransistorNmos: 5.38281e+07 muA
** NormalTransistorNmos: 5.38281e+07 muA
** NormalTransistorNmos: 7.68631e+07 muA
** DiodeTransistorNmos: 7.68621e+07 muA
** NormalTransistorNmos: 3.84321e+07 muA
** NormalTransistorNmos: 3.84321e+07 muA
** NormalTransistorNmos: 8.83346e+08 muA
** NormalTransistorNmos: 8.83345e+08 muA
** NormalTransistorPmos: -8.83345e+08 muA
** DiodeTransistorNmos: 2.10886e+08 muA
** NormalTransistorNmos: 2.10885e+08 muA
** DiodeTransistorNmos: 6.04794e+08 muA
** DiodeTransistorNmos: 2.54483e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.20001  V
** outSourceVoltageBiasXXnXX1: 0.600001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 1.06301  V
** outVoltageBiasXXnXX3: 0.570001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.20801  V
** sourceGCC2: 4.20801  V
** sourceTransconductance: 1.41801  V
** innerStageBias: 0.374001  V
** inner: 0.600001  V


.END