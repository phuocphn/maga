** Name: two_stage_single_output_op_amp_37_12

.MACRO two_stage_single_output_op_amp_37_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=11e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=36e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=431e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=37e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=169e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=59e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=72e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=36e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=308e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=431e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=59e-6
mMainBias14 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=44e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=96e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=96e-6
mSimpleFirstStageLoad17 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=102e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=450e-6
mMainBias19 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=139e-6
mSecondStage1Transconductor20 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad21 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=102e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14e-12
.EOM two_stage_single_output_op_amp_37_12

** Expected Performance Values: 
** Gain: 141 dB
** Power consumption: 8.86801 mW
** Area: 8969 (mu_m)^2
** Transit frequency: 8.48901 MHz
** Transit frequency with error factor: 8.48487 MHz
** Slew rate: 8.00083 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** negPSRR: 108 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 1.06001 V
** VcmMax: 4.83001 V
** VcmMin: 1.35001 V


** Expected Currents: 
** NormalTransistorNmos: 2.88941e+07 muA
** NormalTransistorNmos: 2.03068e+08 muA
** NormalTransistorPmos: -1.0768e+08 muA
** NormalTransistorPmos: -5.61879e+07 muA
** NormalTransistorPmos: -5.61889e+07 muA
** NormalTransistorPmos: -5.61879e+07 muA
** NormalTransistorPmos: -5.61889e+07 muA
** NormalTransistorNmos: 1.12374e+08 muA
** NormalTransistorNmos: 1.12373e+08 muA
** NormalTransistorNmos: 5.61871e+07 muA
** NormalTransistorNmos: 5.61871e+07 muA
** NormalTransistorNmos: 1.3116e+09 muA
** DiodeTransistorNmos: 1.3116e+09 muA
** NormalTransistorPmos: -1.31159e+09 muA
** NormalTransistorPmos: -1.31159e+09 muA
** DiodeTransistorNmos: 1.07681e+08 muA
** NormalTransistorNmos: 1.0768e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.88949e+07 muA
** DiodeTransistorPmos: -2.03067e+08 muA


** Expected Voltages: 
** ibias: 1.14201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.46401  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.03401  V
** outSourceVoltageBiasXXnXX1: 0.732001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX0: 3.96901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.501001  V
** innerTransistorStack1Load1: 4.42501  V
** innerTransistorStack2Load1: 4.42501  V
** out1: 3.86501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.59801  V
** inner: 0.732001  V


.END