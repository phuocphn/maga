** Name: two_stage_single_output_op_amp_114_11

.MACRO two_stage_single_output_op_amp_114_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=2e-6 W=8e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=311e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=92e-6
mTelescopicFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=149e-6
mMainBias5 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=47e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSecondStage1StageBias8 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mTelescopicFirstStageLoad9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=9e-6 W=45e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=10e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=326e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=92e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=23e-6
mMainBias15 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=341e-6
mSecondStage1StageBias16 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=338e-6
mTelescopicFirstStageLoad17 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=9e-6 W=45e-6
mTelescopicFirstStageStageBias18 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=149e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=359e-6
mMainBias20 inputVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=46e-6
mSecondStage1Transconductor21 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad22 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=47e-6
mMainBias23 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=30e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.60001e-12
.EOM two_stage_single_output_op_amp_114_11

** Expected Performance Values: 
** Gain: 149 dB
** Power consumption: 5.76201 mW
** Area: 8490 (mu_m)^2
** Transit frequency: 2.65101 MHz
** Transit frequency with error factor: 2.65013 MHz
** Slew rate: 11.5466 V/mu_s
** Phase margin: 60.1606°
** CMRR: 82 dB
** VoutMax: 4.53001 V
** VoutMin: 0.710001 V
** VcmMax: 4.48001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 2.30181e+07 muA
** NormalTransistorNmos: 3.38446e+08 muA
** NormalTransistorPmos: -1.75226e+08 muA
** NormalTransistorPmos: -2.64741e+08 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 9.52401e+06 muA
** DiodeTransistorPmos: -9.52499e+06 muA
** NormalTransistorPmos: -9.52499e+06 muA
** NormalTransistorNmos: 2.83791e+08 muA
** DiodeTransistorNmos: 2.83791e+08 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 3.21883e+08 muA
** NormalTransistorNmos: 3.21882e+08 muA
** NormalTransistorPmos: -3.21882e+08 muA
** NormalTransistorPmos: -3.21883e+08 muA
** DiodeTransistorNmos: 1.75227e+08 muA
** NormalTransistorNmos: 1.75227e+08 muA
** DiodeTransistorNmos: 2.64742e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.30189e+07 muA
** DiodeTransistorPmos: -3.38445e+08 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 2.65001  V
** inputVoltageBiasXXpXX0: 3.29601  V
** inputVoltageBiasXXpXX1: 1.93601  V
** out: 2.5  V
** outFirstStage: 4.21101  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX3: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.22201  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.579001  V
** innerTransconductance: 2.74401  V
** inner: 0.555001  V


.END