** Name: two_stage_single_output_op_amp_20_6

.MACRO two_stage_single_output_op_amp_20_6 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=119e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=24e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mMainBias4 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=1e-6 W=10e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=156e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=520e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=594e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=119e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=315e-6
mSecondStage1Transconductor10 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=528e-6
mSimpleFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=79e-6
mMainBias12 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=18e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=99e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=520e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=156e-6
mMainBias16 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias17 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=594e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=99e-6
mMainBias19 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=90e-6
mMainBias20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.90001e-12
.EOM two_stage_single_output_op_amp_20_6

** Expected Performance Values: 
** Gain: 142 dB
** Power consumption: 5.25901 mW
** Area: 6974 (mu_m)^2
** Transit frequency: 10.3511 MHz
** Transit frequency with error factor: 10.3365 MHz
** Slew rate: 21.3945 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** negPSRR: 95 dB
** posPSRR: 102 dB
** VoutMax: 3.96001 V
** VoutMin: 0.380001 V
** VcmMax: 3.12001 V
** VcmMin: 0.25 V


** Expected Currents: 
** NormalTransistorNmos: 6.85261e+07 muA
** NormalTransistorPmos: -9.12489e+07 muA
** NormalTransistorPmos: -4.31209e+07 muA
** DiodeTransistorNmos: 1.13327e+08 muA
** NormalTransistorNmos: 1.13327e+08 muA
** NormalTransistorNmos: 1.13327e+08 muA
** NormalTransistorPmos: -2.26654e+08 muA
** DiodeTransistorPmos: -2.26655e+08 muA
** NormalTransistorPmos: -1.13326e+08 muA
** NormalTransistorPmos: -1.13326e+08 muA
** NormalTransistorNmos: 6.02244e+08 muA
** NormalTransistorNmos: 6.02243e+08 muA
** NormalTransistorPmos: -6.02243e+08 muA
** DiodeTransistorPmos: -6.02242e+08 muA
** DiodeTransistorNmos: 9.12481e+07 muA
** DiodeTransistorNmos: 4.31201e+07 muA
** DiodeTransistorPmos: -6.85269e+07 muA
** NormalTransistorPmos: -6.85269e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.56001  V
** outSourceVoltageBiasXXpXX1: 4.28001  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 1.07301  V
** outVoltageBiasXXnXX1: 0.815001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.50101  V
** innerTransconductance: 0.177001  V
** inner: 4.28001  V
** inner: 4.19601  V


.END