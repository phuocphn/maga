** Name: two_stage_single_output_op_amp_31_10

.MACRO two_stage_single_output_op_amp_31_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=6e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=99e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=5e-6 W=380e-6
mMainBias4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSecondStage1StageBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=58e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=54e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=141e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=231e-6
mMainBias9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=16e-6
mMainBias10 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=358e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=599e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=141e-6
mSimpleFirstStageLoad13 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=5e-6 W=380e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=581e-6
mSecondStage1Transconductor15 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=552e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=81e-6
mMainBias17 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=176e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.2001e-12
.EOM two_stage_single_output_op_amp_31_10

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 9.50401 mW
** Area: 14976 (mu_m)^2
** Transit frequency: 5.20201 MHz
** Transit frequency with error factor: 5.19912 MHz
** Slew rate: 4.90248 V/mu_s
** Phase margin: 60.1606°
** CMRR: 108 dB
** negPSRR: 111 dB
** posPSRR: 102 dB
** VoutMax: 4.25 V
** VoutMin: 0.280001 V
** VcmMax: 4.48001 V
** VcmMin: 1.45001 V


** Expected Currents: 
** NormalTransistorNmos: 2.67831e+07 muA
** NormalTransistorNmos: 5.88897e+08 muA
** NormalTransistorPmos: -2.01667e+08 muA
** NormalTransistorPmos: -4.47599e+07 muA
** NormalTransistorPmos: -4.47599e+07 muA
** DiodeTransistorPmos: -4.47599e+07 muA
** NormalTransistorNmos: 8.95171e+07 muA
** NormalTransistorNmos: 8.95161e+07 muA
** NormalTransistorNmos: 4.47591e+07 muA
** NormalTransistorNmos: 4.47591e+07 muA
** NormalTransistorNmos: 9.83986e+08 muA
** NormalTransistorPmos: -9.83985e+08 muA
** NormalTransistorPmos: -9.83986e+08 muA
** DiodeTransistorNmos: 2.01668e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.67839e+07 muA
** DiodeTransistorPmos: -5.88896e+08 muA


** Expected Voltages: 
** ibias: 0.685001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.18201  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.00101  V
** outVoltageBiasXXnXX1: 0.898001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.280001  V
** innerTransistorStack2Load1: 4.25401  V
** out1: 3.51401  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.56501  V


.END