** Name: two_stage_single_output_op_amp_87_3

.MACRO two_stage_single_output_op_amp_87_3 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=94e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=12e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=89e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=46e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=5e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=94e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=309e-6
mTelescopicFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=157e-6
mMainBias10 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=332e-6
mMainBias11 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=496e-6
mTelescopicFirstStageLoad12 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=33e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=74e-6
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=74e-6
mSecondStage1StageBias15 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=575e-6
mMainBias16 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=17e-6
mSecondStage1StageBias17 out outVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=598e-6
mTelescopicFirstStageLoad18 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=33e-6
mMainBias19 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=65e-6
mTelescopicFirstStageStageBias20 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=348e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.6001e-12
.EOM two_stage_single_output_op_amp_87_3

** Expected Performance Values: 
** Gain: 154 dB
** Power consumption: 3.70501 mW
** Area: 14996 (mu_m)^2
** Transit frequency: 5.94801 MHz
** Transit frequency with error factor: 5.94796 MHz
** Slew rate: 9.84774 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 4.41001 V
** VoutMin: 0.150001 V
** VcmMax: 3.99001 V
** VcmMin: 0.370001 V


** Expected Currents: 
** NormalTransistorNmos: 1.25835e+08 muA
** NormalTransistorNmos: 1.88026e+08 muA
** NormalTransistorPmos: -3.40429e+07 muA
** NormalTransistorPmos: -9.08299e+06 muA
** NormalTransistorPmos: -3.00529e+07 muA
** NormalTransistorPmos: -3.00529e+07 muA
** DiodeTransistorNmos: 3.00521e+07 muA
** NormalTransistorNmos: 3.00521e+07 muA
** NormalTransistorNmos: 3.00521e+07 muA
** NormalTransistorPmos: -1.85941e+08 muA
** NormalTransistorPmos: -3.00539e+07 muA
** NormalTransistorPmos: -3.00539e+07 muA
** NormalTransistorNmos: 3.03882e+08 muA
** NormalTransistorPmos: -3.03881e+08 muA
** NormalTransistorPmos: -3.03882e+08 muA
** DiodeTransistorNmos: 3.40421e+07 muA
** DiodeTransistorNmos: 9.08201e+06 muA
** DiodeTransistorPmos: -1.25834e+08 muA
** DiodeTransistorPmos: -1.88025e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.557001  V
** outVoltageBiasXXnXX0: 0.582001  V
** outVoltageBiasXXpXX1: 2.25701  V
** outVoltageBiasXXpXX2: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21401  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 3.04601  V
** sourceGCC2: 3.04601  V
** innerStageBias: 2.79101  V


.END