** Name: two_stage_single_output_op_amp_58_8

.MACRO two_stage_single_output_op_amp_58_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=23e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=71e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=84e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=17e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=32e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=32e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=186e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=179e-6
mFoldedCascodeFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=50e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=50e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=84e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mMainBias16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=92e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=563e-6
mFoldedCascodeFirstStageLoad18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=71e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_58_8

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 2.71601 mW
** Area: 2520 (mu_m)^2
** Transit frequency: 4.74901 MHz
** Transit frequency with error factor: 4.74115 MHz
** Slew rate: 8.96953 V/mu_s
** Phase margin: 73.3387°
** CMRR: 99 dB
** VoutMax: 4.81001 V
** VoutMin: 0.710001 V
** VcmMax: 3 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -4.38079e+07 muA
** NormalTransistorNmos: 4.05651e+07 muA
** NormalTransistorNmos: 6.09491e+07 muA
** NormalTransistorNmos: 4.05651e+07 muA
** NormalTransistorNmos: 6.09491e+07 muA
** DiodeTransistorPmos: -4.05659e+07 muA
** NormalTransistorPmos: -4.05659e+07 muA
** NormalTransistorPmos: -4.07649e+07 muA
** DiodeTransistorPmos: -4.07639e+07 muA
** NormalTransistorPmos: -2.03829e+07 muA
** NormalTransistorPmos: -2.03829e+07 muA
** NormalTransistorNmos: 3.57412e+08 muA
** NormalTransistorNmos: 3.57411e+08 muA
** NormalTransistorPmos: -3.57411e+08 muA
** DiodeTransistorNmos: 4.38071e+07 muA
** DiodeTransistorNmos: 4.38071e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.30201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11001  V
** out: 2.5  V
** outFirstStage: 4.24701  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.25701  V
** sourceGCC1: 0.537001  V
** sourceGCC2: 0.537001  V
** sourceTransconductance: 3.36501  V
** innerStageBias: 0.551001  V
** inner: 4.14801  V


.END