** Name: two_stage_single_output_op_amp_11_8

.MACRO two_stage_single_output_op_amp_11_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=35e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=14e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=6e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=369e-6
mSecondStage1StageBias9 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=7e-6 W=257e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=6e-6
mMainBias11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=120e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=35e-6
mMainBias15 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=60e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_11_8

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 3.48401 mW
** Area: 3582 (mu_m)^2
** Transit frequency: 2.95301 MHz
** Transit frequency with error factor: 2.94876 MHz
** Slew rate: 7.64592 V/mu_s
** Phase margin: 67.0361°
** CMRR: 97 dB
** negPSRR: 90 dB
** posPSRR: 85 dB
** VoutMax: 4.25 V
** VoutMin: 0.640001 V
** VcmMax: 3.64001 V
** VcmMin: 1.02001 V


** Expected Currents: 
** NormalTransistorNmos: 8.21501e+06 muA
** NormalTransistorPmos: -3.49139e+07 muA
** DiodeTransistorPmos: -1.72509e+07 muA
** DiodeTransistorPmos: -1.72519e+07 muA
** NormalTransistorPmos: -1.72509e+07 muA
** NormalTransistorPmos: -1.72519e+07 muA
** NormalTransistorNmos: 3.45011e+07 muA
** NormalTransistorNmos: 1.72501e+07 muA
** NormalTransistorNmos: 1.72501e+07 muA
** NormalTransistorNmos: 6.09204e+08 muA
** NormalTransistorNmos: 6.09203e+08 muA
** NormalTransistorPmos: -6.09203e+08 muA
** DiodeTransistorNmos: 3.49131e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.21599e+06 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 1.04401  V
** outVoltageBiasXXpXX0: 3.99201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.23801  V
** innerSourceLoad1: 4.03601  V
** innerTransistorStack2Load1: 4.03601  V
** sourceTransconductance: 1.68101  V
** innerStageBias: 0.198001  V


.END