** Name: two_stage_single_output_op_amp_55_12

.MACRO two_stage_single_output_op_amp_55_12 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=97e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=97e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=14e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=71e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=36e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=97e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=195e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=195e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=155e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=71e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=3e-6 W=97e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=482e-6
mMainBias16 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=100e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerOutputLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=227e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=132e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=132e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=443e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=227e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=222e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.2001e-12
.EOM two_stage_single_output_op_amp_55_12

** Expected Performance Values: 
** Gain: 172 dB
** Power consumption: 11.5271 mW
** Area: 9512 (mu_m)^2
** Transit frequency: 6.47101 MHz
** Transit frequency with error factor: 6.47099 MHz
** Slew rate: 5.0409 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 1.71001 V
** VcmMax: 5.15001 V
** VcmMin: 0.75 V


** Expected Currents: 
** NormalTransistorNmos: 3.65522e+08 muA
** NormalTransistorNmos: 7.56941e+07 muA
** NormalTransistorPmos: -2.56004e+08 muA
** NormalTransistorPmos: -9.21919e+07 muA
** NormalTransistorPmos: -1.50813e+08 muA
** NormalTransistorPmos: -9.21919e+07 muA
** NormalTransistorPmos: -1.50813e+08 muA
** DiodeTransistorNmos: 9.21911e+07 muA
** NormalTransistorNmos: 9.21901e+07 muA
** NormalTransistorNmos: 9.21911e+07 muA
** DiodeTransistorNmos: 9.21901e+07 muA
** NormalTransistorNmos: 1.17244e+08 muA
** NormalTransistorNmos: 5.86211e+07 muA
** NormalTransistorNmos: 5.86211e+07 muA
** NormalTransistorNmos: 1.29656e+09 muA
** DiodeTransistorNmos: 1.29656e+09 muA
** NormalTransistorPmos: -1.29655e+09 muA
** NormalTransistorPmos: -1.29656e+09 muA
** DiodeTransistorNmos: 2.56005e+08 muA
** NormalTransistorNmos: 2.56004e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.65521e+08 muA
** DiodeTransistorPmos: -7.56949e+07 muA


** Expected Voltages: 
** ibias: 0.595001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.03201  V
** outInputVoltageBiasXXnXX1: 2.11801  V
** outSourceVoltageBiasXXnXX1: 1.05901  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.18201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.20401  V
** innerSourceLoad2: 0.616001  V
** innerTransistorStack1Load2: 0.615001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.93701  V
** innerTransconductance: 4.59601  V
** inner: 1.05301  V


.END