** Name: two_stage_single_output_op_amp_79_11

.MACRO two_stage_single_output_op_amp_79_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=14e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=39e-6
mFoldedCascodeFirstStageStageBias5 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=27e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=7e-6 W=59e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=40e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=40e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=44e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=359e-6
mSecondStage1StageBias13 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=7e-6 W=583e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=59e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=524e-6
mMainBias16 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=41e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=161e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=161e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=389e-6
mMainBias21 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=152e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=188e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=41e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_79_11

** Expected Performance Values: 
** Gain: 185 dB
** Power consumption: 3.61601 mW
** Area: 13763 (mu_m)^2
** Transit frequency: 4.46901 MHz
** Transit frequency with error factor: 4.46901 MHz
** Slew rate: 3.68017 V/mu_s
** Phase margin: 64.7443°
** CMRR: 146 dB
** VoutMax: 4.54001 V
** VoutMin: 0.350001 V
** VcmMax: 5.13001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 3.75676e+08 muA
** NormalTransistorNmos: 6.40801e+06 muA
** NormalTransistorPmos: -2.51869e+07 muA
** NormalTransistorPmos: -1.66509e+07 muA
** NormalTransistorPmos: -2.61859e+07 muA
** NormalTransistorPmos: -1.66509e+07 muA
** NormalTransistorPmos: -2.61859e+07 muA
** NormalTransistorNmos: 1.66501e+07 muA
** NormalTransistorNmos: 1.66491e+07 muA
** NormalTransistorNmos: 1.66501e+07 muA
** NormalTransistorNmos: 1.66491e+07 muA
** NormalTransistorNmos: 1.90691e+07 muA
** NormalTransistorNmos: 1.90701e+07 muA
** NormalTransistorNmos: 9.53401e+06 muA
** NormalTransistorNmos: 9.53401e+06 muA
** NormalTransistorNmos: 2.53558e+08 muA
** NormalTransistorNmos: 2.53557e+08 muA
** NormalTransistorPmos: -2.53557e+08 muA
** NormalTransistorPmos: -2.53558e+08 muA
** DiodeTransistorNmos: 2.51861e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.75675e+08 muA
** DiodeTransistorPmos: -6.40899e+06 muA


** Expected Voltages: 
** ibias: 0.564001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.953001  V
** out: 2.5  V
** outFirstStage: 4.24501  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.16501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.359001  V
** innerTransistorStack1Load2: 0.395001  V
** innerTransistorStack2Load2: 0.395001  V
** out1: 0.599001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.359001  V
** innerTransconductance: 4.52401  V


.END