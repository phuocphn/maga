** Name: two_stage_single_output_op_amp_6_3

.MACRO two_stage_single_output_op_amp_6_3 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=122e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=4e-6 W=122e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=76e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=112e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=4e-6 W=122e-6
mMainBias7 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=360e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=194e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=122e-6
mSimpleFirstStageTransconductor10 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=79e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=163e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=417e-6
mMainBias13 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=286e-6
mSecondStage1StageBias14 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=598e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=79e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.70001e-12
.EOM two_stage_single_output_op_amp_6_3

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 9.41101 mW
** Area: 9148 (mu_m)^2
** Transit frequency: 4.03901 MHz
** Transit frequency with error factor: 4.02559 MHz
** Slew rate: 12.4011 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** negPSRR: 88 dB
** posPSRR: 93 dB
** VoutMax: 4.52001 V
** VoutMin: 0.330001 V
** VcmMax: 3.44001 V
** VcmMin: 0.570001 V


** Expected Currents: 
** NormalTransistorNmos: 1.13719e+09 muA
** NormalTransistorPmos: -2.41694e+08 muA
** DiodeTransistorNmos: 6.88741e+07 muA
** NormalTransistorNmos: 6.88731e+07 muA
** NormalTransistorNmos: 6.88741e+07 muA
** DiodeTransistorNmos: 6.88731e+07 muA
** NormalTransistorPmos: -1.37748e+08 muA
** NormalTransistorPmos: -6.8875e+07 muA
** NormalTransistorPmos: -6.8875e+07 muA
** NormalTransistorNmos: 3.45601e+08 muA
** NormalTransistorPmos: -3.456e+08 muA
** NormalTransistorPmos: -3.45601e+08 muA
** DiodeTransistorNmos: 2.41695e+08 muA
** DiodeTransistorPmos: -1.13718e+09 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.837001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.731001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 1.13601  V
** innerTransistorStack1Load1: 0.567001  V
** innerTransistorStack2Load1: 0.568001  V
** sourceTransconductance: 3.75901  V
** innerStageBias: 4.42901  V


.END