** Name: two_stage_single_output_op_amp_159_4

.MACRO two_stage_single_output_op_amp_159_4 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=56e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=106e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=544e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=14e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=62e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=162e-6
mSecondStage1Transconductor8 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=71e-6
mSimpleFirstStageLoad9 outFirstStage outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=62e-6
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=104e-6
mSimpleFirstStageLoad12 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=544e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=13e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=306e-6
mMainBias15 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=519e-6
mSecondStage1StageBias16 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=595e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=7e-6 W=128e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=104e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=203e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_159_4

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 6.47301 mW
** Area: 11876 (mu_m)^2
** Transit frequency: 4.06201 MHz
** Transit frequency with error factor: 4.04523 MHz
** Slew rate: 3.9987 V/mu_s
** Phase margin: 67.6091°
** CMRR: 95 dB
** VoutMax: 4.03001 V
** VoutMin: 0.470001 V
** VcmMax: 3.20001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -5.26202e+08 muA
** NormalTransistorPmos: -2.01891e+08 muA
** NormalTransistorPmos: -1.08962e+08 muA
** NormalTransistorPmos: -1.08962e+08 muA
** DiodeTransistorPmos: -1.08962e+08 muA
** NormalTransistorNmos: 1.18088e+08 muA
** NormalTransistorNmos: 1.18088e+08 muA
** NormalTransistorPmos: -1.825e+07 muA
** NormalTransistorPmos: -1.82489e+07 muA
** NormalTransistorPmos: -9.125e+06 muA
** NormalTransistorPmos: -9.125e+06 muA
** NormalTransistorNmos: 3.10247e+08 muA
** NormalTransistorNmos: 3.10246e+08 muA
** NormalTransistorPmos: -3.10246e+08 muA
** NormalTransistorPmos: -3.10245e+08 muA
** DiodeTransistorNmos: 5.26203e+08 muA
** DiodeTransistorNmos: 2.01892e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.43501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.875  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.15501  V
** innerStageBias: 4.27801  V
** out1: 3.01101  V
** sourceTransconductance: 3.22001  V
** innerStageBias: 4.16901  V
** innerTransconductance: 0.150001  V


.END