** Name: two_stage_single_output_op_amp_19_3

.MACRO two_stage_single_output_op_amp_19_3 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=74e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=18e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=74e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=132e-6
mSimpleFirstStageLoad7 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=13e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=119e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=28e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=250e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=600e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=119e-6
mMainBias14 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=66e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_19_3

** Expected Performance Values: 
** Gain: 105 dB
** Power consumption: 1.85901 mW
** Area: 4075 (mu_m)^2
** Transit frequency: 5.24701 MHz
** Transit frequency with error factor: 5.24332 MHz
** Slew rate: 6.94231 V/mu_s
** Phase margin: 70.4739°
** CMRR: 104 dB
** negPSRR: 105 dB
** posPSRR: 156 dB
** VoutMax: 4.05001 V
** VoutMin: 0.150001 V
** VcmMax: 3.18001 V
** VcmMin: 0.260001 V


** Expected Currents: 
** NormalTransistorPmos: -6.69149e+07 muA
** DiodeTransistorNmos: 1.57151e+07 muA
** NormalTransistorNmos: 1.57151e+07 muA
** NormalTransistorNmos: 1.57151e+07 muA
** NormalTransistorPmos: -3.14309e+07 muA
** NormalTransistorPmos: -3.14299e+07 muA
** NormalTransistorPmos: -1.57159e+07 muA
** NormalTransistorPmos: -1.57159e+07 muA
** NormalTransistorNmos: 2.5347e+08 muA
** NormalTransistorPmos: -2.53469e+08 muA
** NormalTransistorPmos: -2.53468e+08 muA
** DiodeTransistorNmos: 6.69141e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.45801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.821001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerStageBias: 4.27201  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.27401  V
** innerStageBias: 4.17501  V


.END