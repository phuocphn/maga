** Name: two_stage_single_output_op_amp_46_9

.MACRO two_stage_single_output_op_amp_46_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=22e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=26e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=569e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=51e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=88e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=23e-6
mMainBias7 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=111e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=34e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=129e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=129e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=22e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=569e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=34e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=88e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=8e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=8e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=7e-6 W=600e-6
mMainBias18 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=346e-6
mMainBias19 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=358e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=80e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=23e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_46_9

** Expected Performance Values: 
** Gain: 112 dB
** Power consumption: 5.27201 mW
** Area: 14994 (mu_m)^2
** Transit frequency: 3.11801 MHz
** Transit frequency with error factor: 3.11773 MHz
** Slew rate: 12.1158 V/mu_s
** Phase margin: 70.4739°
** CMRR: 124 dB
** VoutMax: 4.25 V
** VoutMin: 0.850001 V
** VcmMax: 3.63001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -3.15339e+07 muA
** NormalTransistorPmos: -3.23809e+07 muA
** NormalTransistorNmos: 5.46851e+07 muA
** NormalTransistorNmos: 8.20261e+07 muA
** NormalTransistorNmos: 5.46871e+07 muA
** NormalTransistorNmos: 8.20281e+07 muA
** DiodeTransistorPmos: -5.46859e+07 muA
** DiodeTransistorPmos: -5.46869e+07 muA
** NormalTransistorPmos: -5.46879e+07 muA
** NormalTransistorPmos: -5.46869e+07 muA
** NormalTransistorPmos: -5.46829e+07 muA
** NormalTransistorPmos: -2.73419e+07 muA
** NormalTransistorPmos: -2.73419e+07 muA
** NormalTransistorNmos: 8.06478e+08 muA
** DiodeTransistorNmos: 8.06477e+08 muA
** NormalTransistorPmos: -8.06477e+08 muA
** DiodeTransistorNmos: 3.15331e+07 muA
** NormalTransistorNmos: 3.15321e+07 muA
** DiodeTransistorNmos: 3.23801e+07 muA
** DiodeTransistorNmos: 3.23791e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.25801  V
** inputVoltageBiasXXnXX2: 1.17001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.630001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.24901  V
** innerTransistorStack2Load2: 4.24901  V
** out1: 3.32201  V
** sourceGCC1: 0.526001  V
** sourceGCC2: 0.526001  V
** sourceTransconductance: 3.68001  V
** inner: 0.627001  V


.END