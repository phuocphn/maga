** Name: two_stage_single_output_op_amp_170_6

.MACRO two_stage_single_output_op_amp_170_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=38e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=20e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mMainBias5 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=2e-6 W=6e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=26e-6
mSimpleFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=232e-6
mSecondStage1StageBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=559e-6
mSimpleFirstStageLoad9 FirstStageYinnerOutputLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=156e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=170e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=170e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=495e-6
mSecondStage1Transconductor13 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=390e-6
mSimpleFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=156e-6
mMainBias15 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=36e-6
mSimpleFirstStageTransconductor16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=333e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSimpleFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=232e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mMainBias20 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mMainBias21 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=20e-6
mSecondStage1StageBias22 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=559e-6
mSimpleFirstStageLoad23 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=20e-6
mSimpleFirstStageTransconductor24 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=333e-6
mMainBias25 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.7001e-12
.EOM two_stage_single_output_op_amp_170_6

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 6.38901 mW
** Area: 14932 (mu_m)^2
** Transit frequency: 3.82701 MHz
** Transit frequency with error factor: 3.8254 MHz
** Slew rate: 10.1224 V/mu_s
** Phase margin: 60.1606°
** CMRR: 70 dB
** VoutMax: 3.56001 V
** VoutMin: 0.530001 V
** VcmMax: 3 V
** VcmMin: -0.199999 V


** Expected Currents: 
** NormalTransistorNmos: 2.35441e+07 muA
** NormalTransistorPmos: -3.33729e+07 muA
** NormalTransistorPmos: -2.49949e+07 muA
** DiodeTransistorPmos: -7.37099e+06 muA
** DiodeTransistorPmos: -7.37199e+06 muA
** NormalTransistorPmos: -7.37099e+06 muA
** NormalTransistorPmos: -7.37199e+06 muA
** NormalTransistorNmos: 1.1281e+08 muA
** NormalTransistorNmos: 1.12809e+08 muA
** NormalTransistorNmos: 1.1281e+08 muA
** NormalTransistorNmos: 1.12809e+08 muA
** NormalTransistorPmos: -2.10878e+08 muA
** DiodeTransistorPmos: -2.10879e+08 muA
** NormalTransistorPmos: -1.05438e+08 muA
** NormalTransistorPmos: -1.05438e+08 muA
** NormalTransistorNmos: 9.50278e+08 muA
** NormalTransistorNmos: 9.50277e+08 muA
** NormalTransistorPmos: -9.50277e+08 muA
** DiodeTransistorPmos: -9.50276e+08 muA
** DiodeTransistorNmos: 3.33721e+07 muA
** DiodeTransistorNmos: 2.49941e+07 muA
** DiodeTransistorPmos: -2.35449e+07 muA
** NormalTransistorPmos: -2.35459e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.933001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.42001  V
** outSourceVoltageBiasXXpXX1: 4.21001  V
** outSourceVoltageBiasXXpXX2: 4.00201  V
** outVoltageBiasXXnXX2: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.06401  V
** innerSourceLoad1: 3.87701  V
** innerTransistorStack1Load2: 0.321001  V
** innerTransistorStack2Load1: 3.87601  V
** innerTransistorStack2Load2: 0.321001  V
** sourceTransconductance: 3.48301  V
** innerTransconductance: 0.150001  V
** inner: 4.20801  V
** inner: 3.99401  V


.END