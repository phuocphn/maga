** Name: two_stage_single_output_op_amp_177_1

.MACRO two_stage_single_output_op_amp_177_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=23e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=42e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=6e-6 W=21e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=21e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=24e-6
mSimpleFirstStageLoad7 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=177e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=186e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=186e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=28e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=201e-6
mSimpleFirstStageLoad12 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=177e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=60e-6
mSimpleFirstStageTransconductor14 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=90e-6
mSimpleFirstStageStageBias15 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=29e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=21e-6
mSimpleFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=4e-6 W=148e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=586e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=6e-6 W=21e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=90e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_177_1

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 2.33801 mW
** Area: 14984 (mu_m)^2
** Transit frequency: 2.59301 MHz
** Transit frequency with error factor: 2.5914 MHz
** Slew rate: 3.80012 V/mu_s
** Phase margin: 62.4525°
** CMRR: 100 dB
** VoutMax: 4.55001 V
** VoutMin: 0.350001 V
** VcmMax: 3.03001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 6.66701e+06 muA
** NormalTransistorNmos: 1.44281e+07 muA
** DiodeTransistorPmos: -3.55359e+07 muA
** NormalTransistorPmos: -3.55359e+07 muA
** NormalTransistorPmos: -3.55359e+07 muA
** DiodeTransistorPmos: -3.55359e+07 muA
** NormalTransistorNmos: 4.42821e+07 muA
** NormalTransistorNmos: 4.42831e+07 muA
** NormalTransistorNmos: 4.42821e+07 muA
** NormalTransistorNmos: 4.42831e+07 muA
** NormalTransistorPmos: -1.74949e+07 muA
** NormalTransistorPmos: -1.74959e+07 muA
** NormalTransistorPmos: -8.74699e+06 muA
** NormalTransistorPmos: -8.74699e+06 muA
** NormalTransistorNmos: 3.47887e+08 muA
** NormalTransistorPmos: -3.47886e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -6.66799e+06 muA
** DiodeTransistorPmos: -1.44289e+07 muA


** Expected Voltages: 
** ibias: 1.16201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.82301  V
** out: 2.5  V
** outFirstStage: 0.757001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX2: 3.98801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerSourceLoad1: 3.68601  V
** innerStageBias: 4.54901  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.603001  V
** innerTransistorStack2Load2: 0.603001  V
** sourceTransconductance: 3.29701  V


.END