** Name: two_stage_single_output_op_amp_81_12

.MACRO two_stage_single_output_op_amp_81_12 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=47e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=47e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=17e-6
mMainBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=137e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=149e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=232e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=47e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=58e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=58e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=95e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias15 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=137e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=5e-6 W=47e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=486e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=89e-6
mFoldedCascodeFirstStageLoad19 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=266e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=579e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=579e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=422e-6
mMainBias23 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=420e-6
mSecondStage1Transconductor24 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad25 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=266e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.4001e-12
.EOM two_stage_single_output_op_amp_81_12

** Expected Performance Values: 
** Gain: 173 dB
** Power consumption: 9.98701 mW
** Area: 10169 (mu_m)^2
** Transit frequency: 6.01401 MHz
** Transit frequency with error factor: 6.01346 MHz
** Slew rate: 5.54257 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 4.25 V
** VoutMin: 1.06001 V
** VcmMax: 5.23001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 2.33528e+08 muA
** NormalTransistorNmos: 4.26061e+07 muA
** NormalTransistorPmos: -1.17934e+08 muA
** NormalTransistorPmos: -1.08031e+08 muA
** NormalTransistorPmos: -1.63267e+08 muA
** NormalTransistorPmos: -1.08031e+08 muA
** NormalTransistorPmos: -1.63267e+08 muA
** DiodeTransistorNmos: 1.08032e+08 muA
** NormalTransistorNmos: 1.08031e+08 muA
** NormalTransistorNmos: 1.08032e+08 muA
** DiodeTransistorNmos: 1.08031e+08 muA
** NormalTransistorNmos: 1.1047e+08 muA
** NormalTransistorNmos: 1.1047e+08 muA
** NormalTransistorNmos: 5.52351e+07 muA
** NormalTransistorNmos: 5.52351e+07 muA
** NormalTransistorNmos: 1.26676e+09 muA
** DiodeTransistorNmos: 1.26676e+09 muA
** NormalTransistorPmos: -1.26675e+09 muA
** NormalTransistorPmos: -1.26675e+09 muA
** DiodeTransistorNmos: 1.17935e+08 muA
** NormalTransistorNmos: 1.17936e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.33527e+08 muA
** DiodeTransistorPmos: -4.26069e+07 muA


** Expected Voltages: 
** ibias: 1.12601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.46801  V
** out: 2.5  V
** outFirstStage: 4.02801  V
** outSourceVoltageBiasXXnXX1: 0.734001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.25801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.733001  V
** innerStageBias: 0.486001  V
** innerTransistorStack1Load2: 0.730001  V
** out1: 1.50501  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.59201  V
** inner: 0.735001  V


.END