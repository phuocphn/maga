** Name: two_stage_single_output_op_amp_47_9

.MACRO two_stage_single_output_op_amp_47_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=9e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=7e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=217e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=120e-6
mMainBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=6e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=14e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=217e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=14e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=150e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=111e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=111e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=53e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=53e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=7e-6 W=391e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=194e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=106e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=150e-6
mMainBias23 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=202e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_47_9

** Expected Performance Values: 
** Gain: 117 dB
** Power consumption: 3.54301 mW
** Area: 13805 (mu_m)^2
** Transit frequency: 2.76501 MHz
** Transit frequency with error factor: 2.76457 MHz
** Slew rate: 7.07014 V/mu_s
** Phase margin: 65.3172°
** CMRR: 129 dB
** VoutMax: 4.25 V
** VoutMin: 1.31001 V
** VcmMax: 3.84001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.99991e+07 muA
** NormalTransistorPmos: -1.70639e+07 muA
** NormalTransistorPmos: -1.61899e+07 muA
** NormalTransistorNmos: 3.21251e+07 muA
** NormalTransistorNmos: 4.85681e+07 muA
** NormalTransistorNmos: 3.21251e+07 muA
** NormalTransistorNmos: 4.85681e+07 muA
** NormalTransistorPmos: -3.21259e+07 muA
** NormalTransistorPmos: -3.21269e+07 muA
** NormalTransistorPmos: -3.21259e+07 muA
** NormalTransistorPmos: -3.21269e+07 muA
** NormalTransistorPmos: -3.28889e+07 muA
** NormalTransistorPmos: -1.64439e+07 muA
** NormalTransistorPmos: -1.64439e+07 muA
** NormalTransistorNmos: 5.3813e+08 muA
** DiodeTransistorNmos: 5.38129e+08 muA
** NormalTransistorPmos: -5.38129e+08 muA
** DiodeTransistorNmos: 1.70631e+07 muA
** NormalTransistorNmos: 1.70621e+07 muA
** DiodeTransistorNmos: 1.61891e+07 muA
** DiodeTransistorNmos: 1.61901e+07 muA
** DiodeTransistorPmos: -2e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.16601  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.71201  V
** outSourceVoltageBiasXXnXX1: 0.856001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.07501  V
** innerTransistorStack1Load2: 4.43901  V
** innerTransistorStack2Load2: 4.43901  V
** sourceGCC1: 0.527001  V
** sourceGCC2: 0.527001  V
** sourceTransconductance: 3.47901  V
** inner: 0.856001  V


.END