** Name: two_stage_single_output_op_amp_95_12

.MACRO two_stage_single_output_op_amp_95_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=10e-6 W=26e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=11e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=568e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=41e-6
mTelescopicFirstStageLoad5 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=81e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=47e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=9e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=7e-6
mTelescopicFirstStageLoad9 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=33e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=11e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=11e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mMainBias13 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=49e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=568e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=33e-6
mMainBias16 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=104e-6
mTelescopicFirstStageStageBias17 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=10e-6 W=375e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=47e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=311e-6
mMainBias20 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=12e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=7e-6 W=600e-6
mTelescopicFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=81e-6
mMainBias23 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.6001e-12
.EOM two_stage_single_output_op_amp_95_12

** Expected Performance Values: 
** Gain: 180 dB
** Power consumption: 7.56301 mW
** Area: 14997 (mu_m)^2
** Transit frequency: 4.18101 MHz
** Transit frequency with error factor: 4.18075 MHz
** Slew rate: 13.6342 V/mu_s
** Phase margin: 60.1606°
** CMRR: 144 dB
** VoutMax: 3.61001 V
** VoutMin: 0.970001 V
** VcmMax: 3.73001 V
** VcmMin: 0.770001 V


** Expected Currents: 
** NormalTransistorNmos: 1.89091e+07 muA
** NormalTransistorNmos: 4.03441e+07 muA
** NormalTransistorPmos: -2.47569e+07 muA
** NormalTransistorPmos: -1.03089e+08 muA
** NormalTransistorNmos: 2.09521e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** DiodeTransistorPmos: -2.09529e+07 muA
** DiodeTransistorPmos: -2.09529e+07 muA
** NormalTransistorPmos: -2.09519e+07 muA
** NormalTransistorPmos: -2.09529e+07 muA
** NormalTransistorNmos: 1.44991e+08 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 1.27364e+09 muA
** DiodeTransistorNmos: 1.27364e+09 muA
** NormalTransistorPmos: -1.27363e+09 muA
** NormalTransistorPmos: -1.27364e+09 muA
** DiodeTransistorNmos: 2.47561e+07 muA
** NormalTransistorNmos: 2.47551e+07 muA
** DiodeTransistorNmos: 1.0309e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.89099e+07 muA
** DiodeTransistorPmos: -4.03449e+07 muA


** Expected Voltages: 
** ibias: 0.618001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.37201  V
** inputVoltageBiasXXpXX0: 3.47101  V
** out: 2.5  V
** outFirstStage: 3.95501  V
** outSourceVoltageBiasXXnXX1: 0.686001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX1: 2.92601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerOutputLoad2: 3.47801  V
** innerTransistorStack1Load2: 4.21201  V
** innerTransistorStack2Load2: 4.21201  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.39801  V
** inner: 0.684001  V


.END