** Name: two_stage_single_output_op_amp_178_4

.MACRO two_stage_single_output_op_amp_178_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=34e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=64e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=64e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=31e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=17e-6
mSimpleFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=94e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSimpleFirstStageLoad9 FirstStageYinnerOutputLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=409e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=272e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=272e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=160e-6
mSecondStage1Transconductor13 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=484e-6
mSimpleFirstStageLoad14 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=409e-6
mMainBias15 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=20e-6
mSimpleFirstStageTransconductor16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=403e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=64e-6
mSimpleFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=94e-6
mSecondStage1StageBias19 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=151e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mMainBias21 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=16e-6
mSecondStage1StageBias22 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=597e-6
mSimpleFirstStageLoad23 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=64e-6
mSimpleFirstStageTransconductor24 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=403e-6
mMainBias25 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.5e-12
.EOM two_stage_single_output_op_amp_178_4

** Expected Performance Values: 
** Gain: 147 dB
** Power consumption: 4.54201 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 3.47901 MHz
** Transit frequency with error factor: 3.47628 MHz
** Slew rate: 5.59821 V/mu_s
** Phase margin: 60.1606°
** CMRR: 100 dB
** VoutMax: 3.72001 V
** VoutMin: 0.300001 V
** VcmMax: 3.12001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorPmos: -1.01809e+07 muA
** NormalTransistorPmos: -3.23799e+07 muA
** DiodeTransistorPmos: -2.07185e+08 muA
** NormalTransistorPmos: -2.07186e+08 muA
** NormalTransistorPmos: -2.07185e+08 muA
** DiodeTransistorPmos: -2.07186e+08 muA
** NormalTransistorNmos: 2.59665e+08 muA
** NormalTransistorNmos: 2.59664e+08 muA
** NormalTransistorNmos: 2.59665e+08 muA
** NormalTransistorNmos: 2.59664e+08 muA
** NormalTransistorPmos: -1.04958e+08 muA
** DiodeTransistorPmos: -1.04959e+08 muA
** NormalTransistorPmos: -5.24789e+07 muA
** NormalTransistorPmos: -5.24789e+07 muA
** NormalTransistorNmos: 3.07485e+08 muA
** NormalTransistorNmos: 3.07484e+08 muA
** NormalTransistorPmos: -3.07484e+08 muA
** NormalTransistorPmos: -3.07483e+08 muA
** DiodeTransistorNmos: 1.01801e+07 muA
** DiodeTransistorNmos: 3.23791e+07 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90489e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.20701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.37001  V
** outSourceVoltageBiasXXpXX1: 4.18501  V
** outSourceVoltageBiasXXpXX2: 3.96101  V
** outVoltageBiasXXnXX1: 0.705001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.52801  V
** innerTransistorStack1Load1: 3.82601  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load1: 3.83201  V
** innerTransistorStack2Load2: 0.150001  V
** sourceTransconductance: 3.31901  V
** innerStageBias: 4.01001  V
** innerTransconductance: 0.150001  V
** inner: 4.18401  V


.END