** Name: two_stage_single_output_op_amp_205_9

.MACRO two_stage_single_output_op_amp_205_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=8e-6 W=10e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=13e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=5e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=200e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=60e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=10e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=24e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=11e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=200e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=8e-6 W=10e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=24e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=50e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=50e-6
mSimpleFirstStageLoad19 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=600e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=25e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=214e-6
mSimpleFirstStageLoad22 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=600e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=27e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.5e-12
.EOM two_stage_single_output_op_amp_205_9

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 6.29901 mW
** Area: 10189 (mu_m)^2
** Transit frequency: 4.24701 MHz
** Transit frequency with error factor: 4.24481 MHz
** Slew rate: 4.00227 V/mu_s
** Phase margin: 60.1606°
** CMRR: 108 dB
** VoutMax: 4.25 V
** VoutMin: 1.53001 V
** VcmMax: 4.72001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorPmos: -2.71999e+07 muA
** NormalTransistorPmos: -2.49439e+07 muA
** DiodeTransistorNmos: 3.92381e+07 muA
** NormalTransistorNmos: 3.92391e+07 muA
** NormalTransistorNmos: 3.92401e+07 muA
** DiodeTransistorNmos: 3.92391e+07 muA
** NormalTransistorPmos: -5.06669e+07 muA
** NormalTransistorPmos: -5.06679e+07 muA
** NormalTransistorPmos: -5.06689e+07 muA
** NormalTransistorPmos: -5.06679e+07 muA
** NormalTransistorNmos: 2.28551e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 1.14281e+07 muA
** NormalTransistorNmos: 1.14281e+07 muA
** NormalTransistorNmos: 1.08642e+09 muA
** DiodeTransistorNmos: 1.08642e+09 muA
** NormalTransistorPmos: -1.08641e+09 muA
** DiodeTransistorNmos: 2.71991e+07 muA
** NormalTransistorNmos: 2.71981e+07 muA
** DiodeTransistorNmos: 2.49431e+07 muA
** DiodeTransistorNmos: 2.49421e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.12401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.11001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.93801  V
** outSourceVoltageBiasXXnXX1: 0.969001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.90501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.08901  V
** innerStageBias: 0.548001  V
** innerTransistorStack1Load1: 1.09001  V
** innerTransistorStack1Load2: 3.84101  V
** innerTransistorStack2Load2: 3.84101  V
** out1: 2.10601  V
** sourceTransconductance: 1.94501  V
** inner: 0.964001  V


.END