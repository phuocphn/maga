** Name: two_stage_single_output_op_amp_74_8

.MACRO two_stage_single_output_op_amp_74_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=69e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=13e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=9e-6 W=10e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=69e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=10e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=21e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=278e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=13e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=9e-6 W=165e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=6e-6 W=15e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=55e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=36e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=36e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=10e-6 W=553e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=55e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mMainBias22 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_74_8

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 3.44801 mW
** Area: 11502 (mu_m)^2
** Transit frequency: 2.57001 MHz
** Transit frequency with error factor: 2.57029 MHz
** Slew rate: 4.94226 V/mu_s
** Phase margin: 67.6091°
** CMRR: 132 dB
** VoutMax: 4.25 V
** VoutMin: 1.47001 V
** VcmMax: 5.17001 V
** VcmMin: 1.76001 V


** Expected Currents: 
** NormalTransistorPmos: -1.72349e+07 muA
** NormalTransistorPmos: -1.78919e+07 muA
** NormalTransistorPmos: -2.23369e+07 muA
** NormalTransistorPmos: -3.64989e+07 muA
** NormalTransistorPmos: -2.23369e+07 muA
** NormalTransistorPmos: -3.64989e+07 muA
** NormalTransistorNmos: 2.23361e+07 muA
** NormalTransistorNmos: 2.23361e+07 muA
** DiodeTransistorNmos: 2.23361e+07 muA
** NormalTransistorNmos: 2.83211e+07 muA
** DiodeTransistorNmos: 2.83201e+07 muA
** NormalTransistorNmos: 1.41611e+07 muA
** NormalTransistorNmos: 1.41611e+07 muA
** NormalTransistorNmos: 5.61483e+08 muA
** NormalTransistorNmos: 5.61482e+08 muA
** NormalTransistorPmos: -5.61482e+08 muA
** DiodeTransistorNmos: 1.72341e+07 muA
** NormalTransistorNmos: 1.72331e+07 muA
** DiodeTransistorNmos: 1.78911e+07 muA
** DiodeTransistorNmos: 1.78901e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.37201  V
** outInputVoltageBiasXXnXX2: 1.70601  V
** outSourceVoltageBiasXXnXX1: 0.686001  V
** outSourceVoltageBiasXXnXX2: 0.867001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.568001  V
** out1: 1.29701  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.70601  V
** innerStageBias: 0.697001  V
** inner: 0.686001  V


.END