** Name: one_stage_single_output_op_amp62

.MACRO one_stage_single_output_op_amp62 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=11e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=296e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=22e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=72e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=14e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=64e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=173e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=173e-6
mFoldedCascodeFirstStageLoad10 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=64e-6
mMainBias11 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=35e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=27e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=296e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=178e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=178e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=72e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=22e-6
mFoldedCascodeFirstStageLoad18 out outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=8e-6 W=229e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp62

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 1.38601 mW
** Area: 5902 (mu_m)^2
** Transit frequency: 3.90101 MHz
** Transit frequency with error factor: 3.90052 MHz
** Slew rate: 3.74541 V/mu_s
** Phase margin: 88.2356°
** CMRR: 143 dB
** VoutMax: 4.45001 V
** VoutMin: 0.760001 V
** VcmMax: 3.03001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.31641e+07 muA
** NormalTransistorNmos: 1.77671e+07 muA
** NormalTransistorNmos: 7.51411e+07 muA
** NormalTransistorNmos: 1.13141e+08 muA
** NormalTransistorNmos: 7.51411e+07 muA
** NormalTransistorNmos: 1.13141e+08 muA
** DiodeTransistorPmos: -7.51419e+07 muA
** NormalTransistorPmos: -7.51419e+07 muA
** NormalTransistorPmos: -7.51419e+07 muA
** NormalTransistorPmos: -7.60009e+07 muA
** DiodeTransistorPmos: -7.60019e+07 muA
** NormalTransistorPmos: -3.8e+07 muA
** NormalTransistorPmos: -3.8e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.31649e+07 muA
** NormalTransistorPmos: -2.31659e+07 muA
** DiodeTransistorPmos: -1.77679e+07 muA


** Expected Voltages: 
** ibias: 1.14201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outInputVoltageBiasXXpXX1: 3.18201  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.09101  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.63201  V
** out1: 4.26801  V
** sourceGCC1: 0.532001  V
** sourceGCC2: 0.532001  V
** sourceTransconductance: 3.21801  V
** inner: 4.08801  V


.END