** Name: two_stage_single_output_op_amp_50_11

.MACRO two_stage_single_output_op_amp_50_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=23e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=71e-6
mFoldedCascodeFirstStageTransconductor6 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=69e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=69e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=61e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=6e-6 W=598e-6
mFoldedCascodeFirstStageLoad11 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=23e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=85e-6
mMainBias13 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=26e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=181e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=202e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=202e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=384e-6
mMainBias18 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=102e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=417e-6
mFoldedCascodeFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=181e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.5e-12
.EOM two_stage_single_output_op_amp_50_11

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 7.55001 mW
** Area: 8744 (mu_m)^2
** Transit frequency: 6.34901 MHz
** Transit frequency with error factor: 6.34411 MHz
** Slew rate: 5.42088 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** VoutMax: 4.25 V
** VoutMin: 0.540001 V
** VcmMax: 5.09001 V
** VcmMin: 0.790001 V


** Expected Currents: 
** NormalTransistorNmos: 1.42147e+08 muA
** NormalTransistorNmos: 4.34701e+07 muA
** NormalTransistorPmos: -6.15269e+07 muA
** NormalTransistorPmos: -7.35099e+07 muA
** NormalTransistorPmos: -1.23618e+08 muA
** NormalTransistorPmos: -7.35099e+07 muA
** NormalTransistorPmos: -1.23618e+08 muA
** DiodeTransistorNmos: 7.35091e+07 muA
** NormalTransistorNmos: 7.35091e+07 muA
** NormalTransistorNmos: 1.00217e+08 muA
** NormalTransistorNmos: 5.01081e+07 muA
** NormalTransistorNmos: 5.01081e+07 muA
** NormalTransistorNmos: 1.00565e+09 muA
** NormalTransistorNmos: 1.00565e+09 muA
** NormalTransistorPmos: -1.00564e+09 muA
** NormalTransistorPmos: -1.00564e+09 muA
** DiodeTransistorNmos: 6.15261e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.42146e+08 muA
** DiodeTransistorPmos: -4.34709e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.14701  V
** out: 2.5  V
** outFirstStage: 4.05201  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.11701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.679001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.90901  V
** innerStageBias: 0.398001  V
** innerTransconductance: 4.61601  V


.END