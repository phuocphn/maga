** Name: one_stage_single_output_op_amp122

.MACRO one_stage_single_output_op_amp122 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=11e-6
mTelescopicFirstStageStageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=244e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=105e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=7e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mTelescopicFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=75e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=15e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=15e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mTelescopicFirstStageLoad10 out outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=75e-6
mMainBias11 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mMainBias12 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
mTelescopicFirstStageStageBias13 sourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=244e-6
mTelescopicFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mTelescopicFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mTelescopicFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=49e-6
mTelescopicFirstStageLoad17 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=49e-6
mMainBias18 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=115e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp122

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 1.23201 mW
** Area: 4097 (mu_m)^2
** Transit frequency: 3.02501 MHz
** Transit frequency with error factor: 3.02534 MHz
** Slew rate: 10.8991 V/mu_s
** Phase margin: 85.3708°
** CMRR: 136 dB
** VoutMax: 4.41001 V
** VoutMin: 1.06001 V
** VcmMax: 4.98001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorNmos: 9.86201e+06 muA
** NormalTransistorNmos: 8.21901e+06 muA
** NormalTransistorPmos: -1.61272e+08 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorPmos: -2.85709e+07 muA
** NormalTransistorPmos: -2.85719e+07 muA
** NormalTransistorPmos: -2.85709e+07 muA
** NormalTransistorPmos: -2.85719e+07 muA
** NormalTransistorNmos: 2.18414e+08 muA
** DiodeTransistorNmos: 2.18415e+08 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 1.61273e+08 muA
** DiodeTransistorPmos: -9.86299e+06 muA
** DiodeTransistorPmos: -8.21999e+06 muA


** Expected Voltages: 
** ibias: 1.16701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.584001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 3.69201  V
** outVoltageBiasXXpXX1: 3.84601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.72201  V
** innerTransistorStack2Load2: 4.72201  V
** out1: 4.15901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.582001  V


.END