** Name: two_stage_single_output_op_amp_129_4

.MACRO two_stage_single_output_op_amp_129_4 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=90e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=23e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=112e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=32e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
mSimpleFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=151e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=290e-6
mSecondStage1Transconductor8 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=388e-6
mSimpleFirstStageLoad9 outFirstStage outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=151e-6
mMainBias10 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=341e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=49e-6
mSimpleFirstStageLoad12 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=112e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=216e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=586e-6
mSecondStage1StageBias15 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=459e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=157e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=49e-6
mMainBias18 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=545e-6
mMainBias19 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=70e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.8001e-12
.EOM two_stage_single_output_op_amp_129_4

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 5.06501 mW
** Area: 12322 (mu_m)^2
** Transit frequency: 2.61601 MHz
** Transit frequency with error factor: 2.60539 MHz
** Slew rate: 4.59639 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.59001 V
** VoutMin: 0.300001 V
** VcmMax: 3.89001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.24909e+08 muA
** NormalTransistorPmos: -1.72709e+08 muA
** NormalTransistorPmos: -2.19869e+07 muA
** NormalTransistorPmos: -1.09575e+08 muA
** NormalTransistorPmos: -1.09575e+08 muA
** DiodeTransistorPmos: -1.09575e+08 muA
** NormalTransistorNmos: 1.43801e+08 muA
** NormalTransistorNmos: 1.43801e+08 muA
** NormalTransistorPmos: -6.84499e+07 muA
** NormalTransistorPmos: -3.42249e+07 muA
** NormalTransistorPmos: -3.42249e+07 muA
** NormalTransistorNmos: 1.85701e+08 muA
** NormalTransistorNmos: 1.857e+08 muA
** NormalTransistorPmos: -1.857e+08 muA
** NormalTransistorPmos: -1.85701e+08 muA
** DiodeTransistorNmos: 1.7271e+08 muA
** DiodeTransistorNmos: 2.19861e+07 muA
** DiodeTransistorPmos: -3.24908e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX1: 0.705001  V
** outVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.81401  V
** out1: 3.05201  V
** sourceTransconductance: 3.34301  V
** innerStageBias: 4.40001  V
** innerTransconductance: 0.150001  V


.END