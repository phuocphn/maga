** Name: two_stage_single_output_op_amp_2_5

.MACRO two_stage_single_output_op_amp_2_5 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=59e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=68e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=113e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=24e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=210e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=59e-6
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=255e-6
mSimpleFirstStageLoad8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=7e-6 W=59e-6
mMainBias9 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=103e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=222e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=7e-6 W=359e-6
mMainBias12 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=24e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=210e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=222e-6
mMainBias15 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=406e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_2_5

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 3.16101 mW
** Area: 14684 (mu_m)^2
** Transit frequency: 6.24001 MHz
** Transit frequency with error factor: 6.23494 MHz
** Slew rate: 7.08293 V/mu_s
** Phase margin: 65.8902°
** CMRR: 105 dB
** negPSRR: 100 dB
** posPSRR: 105 dB
** VoutMax: 3 V
** VoutMin: 0.300001 V
** VcmMax: 4.07001 V
** VcmMin: 0.140001 V


** Expected Currents: 
** NormalTransistorNmos: 5.47261e+07 muA
** NormalTransistorPmos: -3.66099e+07 muA
** NormalTransistorNmos: 1.61851e+07 muA
** NormalTransistorNmos: 1.61851e+07 muA
** DiodeTransistorNmos: 1.61851e+07 muA
** NormalTransistorPmos: -3.23709e+07 muA
** NormalTransistorPmos: -1.61859e+07 muA
** NormalTransistorPmos: -1.61859e+07 muA
** NormalTransistorNmos: 4.88537e+08 muA
** NormalTransistorPmos: -4.88536e+08 muA
** DiodeTransistorPmos: -4.88536e+08 muA
** DiodeTransistorNmos: 3.66091e+07 muA
** DiodeTransistorPmos: -5.47269e+07 muA
** NormalTransistorPmos: -5.47279e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outInputVoltageBiasXXpXX1: 2.43601  V
** outSourceVoltageBiasXXpXX1: 3.71801  V
** outVoltageBiasXXnXX0: 0.583001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** out1: 1.11001  V
** sourceTransconductance: 3.24401  V
** inner: 3.71101  V


.END