** Name: two_stage_single_output_op_amp_143_10

.MACRO two_stage_single_output_op_amp_143_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=8e-6 W=31e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=353e-6
mSecondStage1StageBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=10e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=8e-6 W=31e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=22e-6
mMainBias8 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=70e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=273e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=10e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=10e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=121e-6
mSimpleFirstStageLoad13 FirstStageYout1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=509e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=588e-6
mSecondStage1Transconductor15 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=548e-6
mSimpleFirstStageLoad16 outFirstStage inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=509e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_143_10

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 4.71701 mW
** Area: 9620 (mu_m)^2
** Transit frequency: 3.50501 MHz
** Transit frequency with error factor: 3.48414 MHz
** Slew rate: 6.64954 V/mu_s
** Phase margin: 76.7764°
** CMRR: 87 dB
** VoutMax: 4.61001 V
** VoutMin: 0.180001 V
** VcmMax: 5.13001 V
** VcmMin: 0.890001 V


** Expected Currents: 
** NormalTransistorNmos: 1.72607e+08 muA
** NormalTransistorNmos: 9.82381e+07 muA
** NormalTransistorNmos: 1.2429e+08 muA
** NormalTransistorNmos: 1.24291e+08 muA
** DiodeTransistorNmos: 1.2429e+08 muA
** NormalTransistorPmos: -1.39726e+08 muA
** NormalTransistorPmos: -1.39726e+08 muA
** NormalTransistorNmos: 3.08751e+07 muA
** NormalTransistorNmos: 1.54371e+07 muA
** NormalTransistorNmos: 1.54371e+07 muA
** NormalTransistorNmos: 3.83126e+08 muA
** NormalTransistorPmos: -3.83125e+08 muA
** NormalTransistorPmos: -3.83126e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.72606e+08 muA
** DiodeTransistorPmos: -9.82389e+07 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.15801  V
** out: 2.5  V
** outFirstStage: 4.24501  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 1.02301  V
** out1: 2.09501  V
** sourceTransconductance: 1.79201  V
** innerTransconductance: 4.44701  V


.END