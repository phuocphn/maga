** Name: two_stage_single_output_op_amp_197_7

.MACRO two_stage_single_output_op_amp_197_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=12e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=19e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias4 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=54e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=11e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=12e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=34e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=5e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=564e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=19e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=34e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=138e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=138e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=402e-6
mMainBias17 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=23e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=360e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=402e-6
mMainBias20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=39e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_197_7

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 7.73601 mW
** Area: 8387 (mu_m)^2
** Transit frequency: 5.92401 MHz
** Transit frequency with error factor: 5.92017 MHz
** Slew rate: 5.58271 V/mu_s
** Phase margin: 61.8795°
** CMRR: 116 dB
** VoutMax: 4.25 V
** VoutMin: 0.160001 V
** VcmMax: 4.60001 V
** VcmMin: 1.61001 V


** Expected Currents: 
** NormalTransistorPmos: -3.60479e+07 muA
** NormalTransistorPmos: -2.11899e+07 muA
** DiodeTransistorNmos: 1.12845e+08 muA
** DiodeTransistorNmos: 1.12846e+08 muA
** NormalTransistorNmos: 1.12845e+08 muA
** NormalTransistorNmos: 1.12846e+08 muA
** NormalTransistorPmos: -1.25796e+08 muA
** NormalTransistorPmos: -1.25797e+08 muA
** NormalTransistorPmos: -1.25796e+08 muA
** NormalTransistorPmos: -1.25797e+08 muA
** NormalTransistorNmos: 2.59031e+07 muA
** NormalTransistorNmos: 2.59021e+07 muA
** NormalTransistorNmos: 1.29521e+07 muA
** NormalTransistorNmos: 1.29521e+07 muA
** NormalTransistorNmos: 1.21841e+09 muA
** NormalTransistorPmos: -1.2184e+09 muA
** DiodeTransistorNmos: 3.60471e+07 muA
** DiodeTransistorNmos: 2.11891e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.564001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 3.93001  V
** outVoltageBiasXXnXX1: 1.05701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15401  V
** innerStageBias: 0.159001  V
** innerTransistorStack1Load2: 3.99701  V
** innerTransistorStack2Load1: 1.15401  V
** innerTransistorStack2Load2: 3.99701  V
** out1: 2.15401  V
** sourceTransconductance: 1.94501  V


.END