** Name: symmetrical_op_amp55

.MACRO symmetrical_op_amp55 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=24e-6
mSecondStage1StageBias5 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=226e-6
mSymmetricalFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=80e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=26e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=26e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=3e-6 W=5e-6
mSecondStage1Transconductor10 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=5e-6
mSymmetricalFirstStageStageBias11 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=80e-6
mMainBias12 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=24e-6
mMainBias13 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=171e-6
mSymmetricalFirstStageTransconductor14 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=125e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias15 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=226e-6
mSecondStage1StageBias16 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=5e-6 W=38e-6
mSymmetricalFirstStageTransconductor17 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=125e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp55

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 1.02401 mW
** Area: 4078 (mu_m)^2
** Transit frequency: 4.21801 MHz
** Transit frequency with error factor: 4.21803 MHz
** Slew rate: 3.93145 V/mu_s
** Phase margin: 85.9437°
** CMRR: 142 dB
** negPSRR: 46 dB
** posPSRR: 48 dB
** VoutMax: 3.70001 V
** VoutMin: 0.720001 V
** VcmMax: 3.19001 V
** VcmMin: 0.0300001 V


** Expected Currents: 
** NormalTransistorPmos: -7.22529e+07 muA
** DiodeTransistorNmos: 1.69001e+07 muA
** DiodeTransistorNmos: 1.69001e+07 muA
** NormalTransistorPmos: -3.38029e+07 muA
** DiodeTransistorPmos: -3.38019e+07 muA
** NormalTransistorPmos: -1.69009e+07 muA
** NormalTransistorPmos: -1.69009e+07 muA
** NormalTransistorNmos: 3.93321e+07 muA
** NormalTransistorNmos: 3.93331e+07 muA
** NormalTransistorPmos: -3.93329e+07 muA
** DiodeTransistorPmos: -3.93339e+07 muA
** NormalTransistorPmos: -3.93349e+07 muA
** NormalTransistorNmos: 3.93341e+07 muA
** NormalTransistorNmos: 3.93331e+07 muA
** DiodeTransistorNmos: 7.22521e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.34001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 1.12101  V
** inSourceTransconductanceComplementarySecondStage: 0.595001  V
** inStageBiasComplementarySecondStage: 4.23801  V
** innerComplementarySecondStage: 3.13401  V
** out: 2.5  V
** outFirstStage: 0.595001  V
** outSourceVoltageBiasXXpXX1: 4.17101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21401  V
** innerTransconductance: 0.190001  V
** inner: 0.190001  V
** inner: 4.16801  V


.END