** Name: two_stage_single_output_op_amp_65_7

.MACRO two_stage_single_output_op_amp_65_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=8e-6 W=155e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=49e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
mMainBias8 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=63e-6
mSecondStage1StageBias9 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=254e-6
mFoldedCascodeFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=49e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=8e-6 W=600e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=133e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=133e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=42e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=42e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=25e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=107e-6
mFoldedCascodeFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=14e-6
mMainBias20 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=368e-6
mMainBias21 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=440e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.10001e-12
.EOM two_stage_single_output_op_amp_65_7

** Expected Performance Values: 
** Gain: 114 dB
** Power consumption: 3.85701 mW
** Area: 14982 (mu_m)^2
** Transit frequency: 2.57601 MHz
** Transit frequency with error factor: 2.57576 MHz
** Slew rate: 4.58882 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 4.29001 V
** VoutMin: 0.150001 V
** VcmMax: 3.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.19993e+08 muA
** NormalTransistorPmos: -2.38119e+07 muA
** NormalTransistorPmos: -2.85709e+07 muA
** NormalTransistorNmos: 2.80521e+07 muA
** NormalTransistorNmos: 4.76161e+07 muA
** NormalTransistorNmos: 2.80521e+07 muA
** NormalTransistorNmos: 4.76161e+07 muA
** NormalTransistorPmos: -2.80529e+07 muA
** NormalTransistorPmos: -2.80539e+07 muA
** NormalTransistorPmos: -2.80529e+07 muA
** NormalTransistorPmos: -2.80539e+07 muA
** NormalTransistorPmos: -3.9125e+07 muA
** NormalTransistorPmos: -3.91239e+07 muA
** NormalTransistorPmos: -1.95629e+07 muA
** NormalTransistorPmos: -1.95629e+07 muA
** NormalTransistorNmos: 4.83776e+08 muA
** NormalTransistorPmos: -4.83775e+08 muA
** DiodeTransistorNmos: 2.38111e+07 muA
** DiodeTransistorNmos: 2.85701e+07 muA
** DiodeTransistorPmos: -1.19992e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.72201  V
** outVoltageBiasXXnXX1: 0.938001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.54501  V
** innerTransistorStack1Load2: 4.58401  V
** innerTransistorStack2Load2: 4.58401  V
** out1: 4.24701  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.45801  V


.END