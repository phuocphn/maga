** Name: two_stage_single_output_op_amp_203_12

.MACRO two_stage_single_output_op_amp_203_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=15e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=15e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=12e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=375e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mSecondStage1StageBias7 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=29e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=330e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=56e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=80e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mMainBias14 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=316e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=375e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=2e-6 W=15e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=56e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=56e-6
mSimpleFirstStageLoad19 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=385e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=377e-6
mSecondStage1Transconductor21 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=385e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=62e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.3001e-12
.EOM two_stage_single_output_op_amp_203_12

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 9.06701 mW
** Area: 14795 (mu_m)^2
** Transit frequency: 5.82901 MHz
** Transit frequency with error factor: 5.81198 MHz
** Slew rate: 5.4936 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** VoutMax: 4.25 V
** VoutMin: 0.950001 V
** VcmMax: 4.88001 V
** VcmMin: 1.42001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorNmos: 1.78961e+07 muA
** NormalTransistorPmos: -3.79579e+07 muA
** DiodeTransistorNmos: 1.79917e+08 muA
** NormalTransistorNmos: 1.79918e+08 muA
** NormalTransistorNmos: 1.79919e+08 muA
** DiodeTransistorNmos: 1.79918e+08 muA
** NormalTransistorPmos: -2.33246e+08 muA
** NormalTransistorPmos: -2.33246e+08 muA
** NormalTransistorNmos: 1.0666e+08 muA
** NormalTransistorNmos: 1.06659e+08 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 1.17942e+09 muA
** DiodeTransistorNmos: 1.17942e+09 muA
** NormalTransistorPmos: -1.17941e+09 muA
** NormalTransistorPmos: -1.17941e+09 muA
** DiodeTransistorNmos: 3.79571e+07 muA
** NormalTransistorNmos: 3.79561e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -1.78969e+07 muA


** Expected Voltages: 
** ibias: 1.17801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.01601  V
** outInputVoltageBiasXXnXX1: 1.35401  V
** outSourceVoltageBiasXXnXX1: 0.677001  V
** outSourceVoltageBiasXXnXX2: 0.556001  V
** outVoltageBiasXXpXX2: 3.91301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.465001  V
** innerTransistorStack1Load1: 1.15601  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.58001  V
** inner: 0.675001  V


.END