** Name: two_stage_single_output_op_amp_152_12

.MACRO two_stage_single_output_op_amp_152_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=7e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=19e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=8e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=132e-6
mMainBias6 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=18e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=300e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=217e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mMainBias12 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=41e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=132e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=7e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=300e-6
mMainBias16 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=502e-6
mSimpleFirstStageLoad17 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=128e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=102e-6
mSimpleFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=102e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=488e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=128e-6
mMainBias23 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=69e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.9001e-12
.EOM two_stage_single_output_op_amp_152_12

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 9.88301 mW
** Area: 14939 (mu_m)^2
** Transit frequency: 6.37801 MHz
** Transit frequency with error factor: 6.37555 MHz
** Slew rate: 6.01127 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** VoutMax: 4.25 V
** VoutMin: 1.61001 V
** VcmMax: 4.66001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorNmos: 2.63988e+08 muA
** NormalTransistorNmos: 2.12391e+07 muA
** NormalTransistorPmos: -8.23599e+07 muA
** DiodeTransistorNmos: 6.37591e+07 muA
** NormalTransistorNmos: 6.37601e+07 muA
** NormalTransistorNmos: 6.37611e+07 muA
** DiodeTransistorNmos: 6.37601e+07 muA
** NormalTransistorPmos: -1.20898e+08 muA
** NormalTransistorPmos: -1.20899e+08 muA
** NormalTransistorPmos: -1.209e+08 muA
** NormalTransistorPmos: -1.20899e+08 muA
** NormalTransistorNmos: 1.14278e+08 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 1.35721e+09 muA
** DiodeTransistorNmos: 1.35721e+09 muA
** NormalTransistorPmos: -1.3572e+09 muA
** NormalTransistorPmos: -1.35721e+09 muA
** DiodeTransistorNmos: 8.23591e+07 muA
** NormalTransistorNmos: 8.23581e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.63987e+08 muA
** DiodeTransistorPmos: -2.12399e+07 muA


** Expected Voltages: 
** ibias: 0.613001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.92001  V
** out: 2.5  V
** outFirstStage: 4.04001  V
** outInputVoltageBiasXXnXX1: 2.01201  V
** outSourceVoltageBiasXXnXX1: 1.00601  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.11801  V
** innerTransistorStack1Load1: 1.14301  V
** innerTransistorStack1Load2: 4.47901  V
** innerTransistorStack2Load1: 1.14201  V
** innerTransistorStack2Load2: 4.47901  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.60401  V
** inner: 1  V


.END