** Name: two_stage_single_output_op_amp_130_5

.MACRO two_stage_single_output_op_amp_130_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=6e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=6e-6 W=22e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=5e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=585e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=11e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=65e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=65e-6
mSimpleFirstStageLoad9 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=67e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=185e-6
mSimpleFirstStageLoad11 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=67e-6
mMainBias12 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mSimpleFirstStageTransconductor14 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=27e-6
mSimpleFirstStageLoad15 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=6e-6 W=22e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=50e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSecondStage1StageBias18 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=585e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=9e-6 W=33e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=27e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_130_5

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 7.13501 mW
** Area: 4559 (mu_m)^2
** Transit frequency: 2.54901 MHz
** Transit frequency with error factor: 2.54752 MHz
** Slew rate: 12.074 V/mu_s
** Phase margin: 73.3387°
** CMRR: 81 dB
** VoutMax: 3.45001 V
** VoutMin: 0.400001 V
** VcmMax: 3.34001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 1.07931e+07 muA
** NormalTransistorNmos: 1.18911e+07 muA
** NormalTransistorPmos: -3.70449e+07 muA
** NormalTransistorPmos: -3.70439e+07 muA
** DiodeTransistorPmos: -3.70449e+07 muA
** NormalTransistorNmos: 6.44581e+07 muA
** NormalTransistorNmos: 6.44571e+07 muA
** NormalTransistorNmos: 6.44571e+07 muA
** NormalTransistorNmos: 6.44571e+07 muA
** NormalTransistorPmos: -5.48289e+07 muA
** NormalTransistorPmos: -2.74139e+07 muA
** NormalTransistorPmos: -2.74139e+07 muA
** NormalTransistorNmos: 1.26535e+09 muA
** NormalTransistorPmos: -1.26534e+09 muA
** DiodeTransistorPmos: -1.26535e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.07939e+07 muA
** NormalTransistorPmos: -1.07949e+07 muA
** DiodeTransistorPmos: -1.18919e+07 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.809001  V
** outInputVoltageBiasXXpXX1: 2.88401  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 3.94201  V
** outVoltageBiasXXpXX2: 4.08701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.605001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.605001  V
** out1: 2.37201  V
** sourceTransconductance: 3.81401  V
** inner: 3.93801  V


.END