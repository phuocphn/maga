** Name: two_stage_single_output_op_amp_189_7

.MACRO two_stage_single_output_op_amp_189_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=53e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=10e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=38e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=457e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=2e-6 W=8e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=38e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=103e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=103e-6
mSimpleFirstStageLoad15 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=67e-6
mMainBias16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=191e-6
mMainBias17 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=84e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=512e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=67e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_189_7

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 6.23801 mW
** Area: 8111 (mu_m)^2
** Transit frequency: 3.76701 MHz
** Transit frequency with error factor: 3.76433 MHz
** Slew rate: 3.5498 V/mu_s
** Phase margin: 65.3172°
** CMRR: 119 dB
** VoutMax: 4.25 V
** VoutMin: 0.340001 V
** VcmMax: 4.87001 V
** VcmMin: 1.49001 V


** Expected Currents: 
** NormalTransistorPmos: -1.92386e+08 muA
** NormalTransistorPmos: -8.45809e+07 muA
** NormalTransistorNmos: 9.59561e+07 muA
** NormalTransistorNmos: 9.59571e+07 muA
** DiodeTransistorNmos: 9.59561e+07 muA
** NormalTransistorPmos: -1.03998e+08 muA
** NormalTransistorPmos: -1.04e+08 muA
** NormalTransistorPmos: -1.04e+08 muA
** NormalTransistorPmos: -1.04e+08 muA
** NormalTransistorNmos: 1.60831e+07 muA
** NormalTransistorNmos: 1.60821e+07 muA
** NormalTransistorNmos: 8.04201e+06 muA
** NormalTransistorNmos: 8.04201e+06 muA
** NormalTransistorNmos: 7.42649e+08 muA
** NormalTransistorPmos: -7.42648e+08 muA
** DiodeTransistorNmos: 1.92387e+08 muA
** DiodeTransistorNmos: 8.45801e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.15501  V
** inputVoltageBiasXXnXX2: 0.743001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.555001  V
** innerTransistorStack1Load2: 4.25601  V
** innerTransistorStack2Load2: 4.25601  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V


.END