** Name: two_stage_single_output_op_amp_72_4

.MACRO two_stage_single_output_op_amp_72_4 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=80e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=289e-6
mFoldedCascodeFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mSecondStage1StageBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=19e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=21e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=40e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=40e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=11e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=97e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=289e-6
mSecondStage1Transconductor12 out outVoltageBiasXXnXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=33e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=80e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=97e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=91e-6
mSecondStage1StageBias18 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=97e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=279e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=132e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_72_4

** Expected Performance Values: 
** Gain: 147 dB
** Power consumption: 5.51701 mW
** Area: 5453 (mu_m)^2
** Transit frequency: 4.28401 MHz
** Transit frequency with error factor: 4.27973 MHz
** Slew rate: 4.14999 V/mu_s
** Phase margin: 60.1606°
** CMRR: 108 dB
** VoutMax: 3.78001 V
** VoutMin: 0.410001 V
** VcmMax: 4.93001 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorPmos: -5.68132e+08 muA
** NormalTransistorPmos: -2.68793e+08 muA
** NormalTransistorPmos: -1.96969e+07 muA
** NormalTransistorPmos: -3.05439e+07 muA
** NormalTransistorPmos: -1.96969e+07 muA
** NormalTransistorPmos: -3.05439e+07 muA
** DiodeTransistorNmos: 1.96961e+07 muA
** NormalTransistorNmos: 1.96961e+07 muA
** NormalTransistorNmos: 2.16911e+07 muA
** DiodeTransistorNmos: 2.16901e+07 muA
** NormalTransistorNmos: 1.08461e+07 muA
** NormalTransistorNmos: 1.08461e+07 muA
** NormalTransistorNmos: 1.85306e+08 muA
** NormalTransistorNmos: 1.85305e+08 muA
** NormalTransistorPmos: -1.85305e+08 muA
** NormalTransistorPmos: -1.85304e+08 muA
** DiodeTransistorNmos: 5.68133e+08 muA
** NormalTransistorNmos: 5.68132e+08 muA
** DiodeTransistorNmos: 2.68794e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.16601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXnXX1: 1.11401  V
** outSourceVoltageBiasXXnXX1: 0.557001  V
** outSourceVoltageBiasXXpXX1: 3.96101  V
** outVoltageBiasXXnXX2: 0.812001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.557001  V
** sourceGCC1: 3.88001  V
** sourceGCC2: 3.88001  V
** sourceTransconductance: 1.92501  V
** innerStageBias: 3.91501  V
** innerTransconductance: 0.150001  V
** inner: 0.556001  V


.END