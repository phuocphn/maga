** Name: two_stage_single_output_op_amp_206_10

.MACRO two_stage_single_output_op_amp_206_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=13e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=13e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=14e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=95e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=34e-6
mMainBias6 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=472e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=69e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=27e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=13e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=34e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=95e-6
mMainBias12 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=471e-6
mSecondStage1StageBias13 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=550e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=1e-6 W=13e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=27e-6
mMainBias16 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=498e-6
mSimpleFirstStageLoad17 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=431e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=470e-6
mSimpleFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=470e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=317e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=252e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=431e-6
mMainBias23 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=102e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_206_10

** Expected Performance Values: 
** Gain: 103 dB
** Power consumption: 9.00101 mW
** Area: 14941 (mu_m)^2
** Transit frequency: 5.87701 MHz
** Transit frequency with error factor: 5.87267 MHz
** Slew rate: 5.53875 V/mu_s
** Phase margin: 60.1606°
** CMRR: 124 dB
** VoutMax: 4.33001 V
** VoutMin: 0.180001 V
** VcmMax: 4.77001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 3.50292e+08 muA
** NormalTransistorNmos: 3.32171e+08 muA
** NormalTransistorPmos: -7.17819e+07 muA
** DiodeTransistorNmos: 3.11857e+08 muA
** NormalTransistorNmos: 3.11858e+08 muA
** NormalTransistorNmos: 3.11859e+08 muA
** DiodeTransistorNmos: 3.11858e+08 muA
** NormalTransistorPmos: -3.24713e+08 muA
** NormalTransistorPmos: -3.24714e+08 muA
** NormalTransistorPmos: -3.24715e+08 muA
** NormalTransistorPmos: -3.24714e+08 muA
** NormalTransistorNmos: 2.57131e+07 muA
** DiodeTransistorNmos: 2.57121e+07 muA
** NormalTransistorNmos: 1.28571e+07 muA
** NormalTransistorNmos: 1.28571e+07 muA
** NormalTransistorNmos: 3.8654e+08 muA
** NormalTransistorPmos: -3.86539e+08 muA
** NormalTransistorPmos: -3.8654e+08 muA
** DiodeTransistorNmos: 7.17811e+07 muA
** NormalTransistorNmos: 7.17801e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.50291e+08 muA
** DiodeTransistorPmos: -3.3217e+08 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.09401  V
** out: 2.5  V
** outFirstStage: 4.17401  V
** outInputVoltageBiasXXnXX1: 1.23201  V
** outSourceVoltageBiasXXnXX1: 0.616001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack1Load1: 1.15601  V
** innerTransistorStack1Load2: 4.53901  V
** innerTransistorStack2Load2: 4.53901  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.66301  V
** inner: 0.615001  V


.END