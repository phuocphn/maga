** Name: symmetrical_op_amp93

.MACRO symmetrical_op_amp93 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=160e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=40e-6
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=40e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=97e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=97e-6
mSymmetricalFirstStageLoad10 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=121e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 inStageBiasComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=3e-6 W=156e-6
mSecondStage1Transconductor12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=156e-6
mSymmetricalFirstStageLoad13 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=121e-6
mMainBias14 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=48e-6
mSymmetricalFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=559e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=160e-6
mSymmetricalFirstStageTransconductor17 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=394e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=68e-6
mSymmetricalFirstStageTransconductor19 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=394e-6
mMainBias20 out2FirstStage ibias sourcePmos sourcePmos pmos4 L=4e-6 W=51e-6
mMainBias21 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=38e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp93

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 3.34701 mW
** Area: 9238 (mu_m)^2
** Transit frequency: 12.6741 MHz
** Transit frequency with error factor: 12.6737 MHz
** Slew rate: 18.43 V/mu_s
** Phase margin: 81.3601°
** CMRR: 145 dB
** negPSRR: 48 dB
** posPSRR: 58 dB
** VoutMax: 4.36001 V
** VoutMin: 0.350001 V
** VcmMax: 3.96001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -1.04609e+07 muA
** NormalTransistorPmos: -1.40219e+07 muA
** NormalTransistorNmos: 7.69481e+07 muA
** NormalTransistorNmos: 7.69471e+07 muA
** NormalTransistorNmos: 7.69481e+07 muA
** NormalTransistorNmos: 7.69471e+07 muA
** NormalTransistorPmos: -1.53897e+08 muA
** NormalTransistorPmos: -7.69489e+07 muA
** NormalTransistorPmos: -7.69489e+07 muA
** NormalTransistorNmos: 1.84749e+08 muA
** NormalTransistorNmos: 1.8475e+08 muA
** NormalTransistorPmos: -1.84748e+08 muA
** NormalTransistorPmos: -1.8475e+08 muA
** DiodeTransistorPmos: -1.84748e+08 muA
** NormalTransistorNmos: 1.84749e+08 muA
** NormalTransistorNmos: 1.8475e+08 muA
** DiodeTransistorNmos: 1.04601e+07 muA
** DiodeTransistorNmos: 1.40211e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18901  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** inStageBiasComplementarySecondStage: 4.18101  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.759001  V
** outVoltageBiasXXnXX0: 0.720001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.204001  V
** innerTransistorStack2Load1: 0.204001  V
** sourceTransconductance: 3.29701  V
** innerStageBias: 4.63801  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END