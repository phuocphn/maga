** Name: two_stage_single_output_op_amp_10_12

.MACRO two_stage_single_output_op_amp_10_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=7e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=141e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=130e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=121e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=19e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mSecondStage1StageBias10 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=141e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=19e-6
mMainBias12 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=210e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=244e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=130e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=570e-6
mSecondStage1Transconductor16 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=583e-6
mSimpleFirstStageLoad17 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=256e-6
mMainBias18 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.4001e-12
.EOM two_stage_single_output_op_amp_10_12

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 8.06101 mW
** Area: 8321 (mu_m)^2
** Transit frequency: 9.34401 MHz
** Transit frequency with error factor: 9.32556 MHz
** Slew rate: 30.7064 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** negPSRR: 114 dB
** posPSRR: 90 dB
** VoutMax: 4.40001 V
** VoutMin: 1.88001 V
** VcmMax: 4.37001 V
** VcmMin: 1.15001 V


** Expected Currents: 
** NormalTransistorNmos: 1.21646e+08 muA
** NormalTransistorNmos: 1.42147e+08 muA
** NormalTransistorPmos: -4.66979e+07 muA
** DiodeTransistorPmos: -1.76713e+08 muA
** NormalTransistorPmos: -1.76713e+08 muA
** NormalTransistorPmos: -1.76713e+08 muA
** NormalTransistorNmos: 3.53426e+08 muA
** NormalTransistorNmos: 1.76714e+08 muA
** NormalTransistorNmos: 1.76714e+08 muA
** NormalTransistorNmos: 9.38379e+08 muA
** DiodeTransistorNmos: 9.38378e+08 muA
** NormalTransistorPmos: -9.38378e+08 muA
** NormalTransistorPmos: -9.38377e+08 muA
** DiodeTransistorNmos: 4.66971e+07 muA
** NormalTransistorNmos: 4.66961e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.21645e+08 muA
** DiodeTransistorPmos: -1.42146e+08 muA


** Expected Voltages: 
** ibias: 0.571001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.13401  V
** outInputVoltageBiasXXnXX1: 2.28801  V
** outSourceVoltageBiasXXnXX1: 1.14401  V
** outVoltageBiasXXpXX0: 4.20001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.15901  V
** innerTransistorStack2Load1: 4.44601  V
** sourceTransconductance: 1.51901  V
** innerTransconductance: 4.54901  V
** inner: 1.13701  V


.END