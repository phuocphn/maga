** Name: two_stage_single_output_op_amp_123_12

.MACRO two_stage_single_output_op_amp_123_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=4e-6 W=14e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=43e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=531e-6
mMainBias4 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=21e-6
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=127e-6
mTelescopicFirstStageLoad7 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=10e-6 W=127e-6
mMainBias8 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=15e-6
mSecondStage1StageBias9 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
mTelescopicFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=412e-6
mTelescopicFirstStageLoad11 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=20e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=20e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=43e-6
mMainBias15 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=18e-6
mSecondStage1StageBias16 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=531e-6
mTelescopicFirstStageLoad17 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
mMainBias18 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=236e-6
mTelescopicFirstStageStageBias19 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=138e-6
mTelescopicFirstStageLoad20 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=127e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=280e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=6e-6 W=542e-6
mTelescopicFirstStageLoad23 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=10e-6 W=127e-6
mMainBias24 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=144e-6
mMainBias25 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=277e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.60001e-12
.EOM two_stage_single_output_op_amp_123_12

** Expected Performance Values: 
** Gain: 180 dB
** Power consumption: 7.10601 mW
** Area: 14983 (mu_m)^2
** Transit frequency: 4.67601 MHz
** Transit frequency with error factor: 4.67645 MHz
** Slew rate: 22.7352 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 3.76001 V
** VoutMin: 0.700001 V
** VcmMax: 3.68001 V
** VcmMin: 1.37001 V


** Expected Currents: 
** NormalTransistorNmos: 8.65701e+06 muA
** NormalTransistorNmos: 1.12815e+08 muA
** NormalTransistorPmos: -8.18999e+07 muA
** NormalTransistorPmos: -1.58405e+08 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90489e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** DiodeTransistorPmos: -1.90489e+07 muA
** NormalTransistorNmos: 1.96499e+08 muA
** NormalTransistorNmos: 1.96498e+08 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.01136e+09 muA
** DiodeTransistorNmos: 1.01136e+09 muA
** NormalTransistorPmos: -1.01135e+09 muA
** NormalTransistorPmos: -1.01135e+09 muA
** DiodeTransistorNmos: 8.18991e+07 muA
** NormalTransistorNmos: 8.18991e+07 muA
** DiodeTransistorNmos: 1.58406e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -8.65799e+06 muA
** DiodeTransistorPmos: -1.12814e+08 muA


** Expected Voltages: 
** ibias: 1.14301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.92901  V
** out: 2.5  V
** outFirstStage: 3.98501  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX3: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX1: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.27701  V
** innerStageBias: 0.478001  V
** innerTransistorStack1Load2: 4.27501  V
** out1: 3.42201  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 3.28801  V
** inner: 0.555001  V


.END