** Name: two_stage_single_output_op_amp_134_6

.MACRO two_stage_single_output_op_amp_134_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=10e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=17e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=17e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=85e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=6e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=126e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=276e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=276e-6
mSimpleFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=72e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=130e-6
mSecondStage1Transconductor12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=8e-6 W=289e-6
mSimpleFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=72e-6
mMainBias14 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=42e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
mSimpleFirstStageTransconductor16 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=33e-6
mSimpleFirstStageStageBias17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=600e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=6e-6
mMainBias19 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=37e-6
mSecondStage1StageBias20 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=126e-6
mSimpleFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=17e-6
mSimpleFirstStageTransconductor22 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=33e-6
mMainBias23 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=475e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7e-12
.EOM two_stage_single_output_op_amp_134_6

** Expected Performance Values: 
** Gain: 134 dB
** Power consumption: 3.63801 mW
** Area: 14992 (mu_m)^2
** Transit frequency: 4.64301 MHz
** Transit frequency with error factor: 4.63867 MHz
** Slew rate: 10.1575 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 3 V
** VoutMin: 0.540001 V
** VcmMax: 3.89001 V
** VcmMin: 0 V


** Expected Currents: 
** NormalTransistorNmos: 1.82921e+07 muA
** NormalTransistorPmos: -5.58539e+07 muA
** NormalTransistorPmos: -4.34599e+06 muA
** DiodeTransistorPmos: -8.63029e+07 muA
** DiodeTransistorPmos: -8.63029e+07 muA
** NormalTransistorPmos: -8.63029e+07 muA
** NormalTransistorPmos: -8.63029e+07 muA
** NormalTransistorNmos: 1.22044e+08 muA
** NormalTransistorNmos: 1.22043e+08 muA
** NormalTransistorNmos: 1.22044e+08 muA
** NormalTransistorNmos: 1.22043e+08 muA
** NormalTransistorPmos: -7.14809e+07 muA
** NormalTransistorPmos: -3.57409e+07 muA
** NormalTransistorPmos: -3.57409e+07 muA
** NormalTransistorNmos: 3.85093e+08 muA
** NormalTransistorNmos: 3.85094e+08 muA
** NormalTransistorPmos: -3.85092e+08 muA
** DiodeTransistorPmos: -3.85093e+08 muA
** DiodeTransistorNmos: 5.58531e+07 muA
** DiodeTransistorNmos: 4.34501e+06 muA
** DiodeTransistorPmos: -1.82929e+07 muA
** NormalTransistorPmos: -1.82939e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.23701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.566001  V
** out: 2.5  V
** outFirstStage: 0.593001  V
** outInputVoltageBiasXXpXX1: 2.43601  V
** outSourceVoltageBiasXXpXX1: 3.71701  V
** outVoltageBiasXXnXX1: 0.965001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.161001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.161001  V
** out1: 2.37201  V
** sourceTransconductance: 3.41101  V
** innerTransconductance: 0.204001  V
** inner: 3.71201  V


.END