** Name: two_stage_single_output_op_amp_76_9

.MACRO two_stage_single_output_op_amp_76_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=43e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=23e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=4e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=30e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=183e-6
mMainBias6 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=36e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=25e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=43e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=30e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=23e-6
mMainBias14 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=183e-6
mFoldedCascodeFirstStageLoad16 outFirstStage outVoltageBiasXXnXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=18e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=221e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=91e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=91e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=369e-6
mFoldedCascodeFirstStageLoad21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=221e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=56e-6
mMainBias23 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=101e-6
mMainBias24 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=596e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_76_9

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 11.3391 mW
** Area: 8626 (mu_m)^2
** Transit frequency: 4.22701 MHz
** Transit frequency with error factor: 4.22701 MHz
** Slew rate: 4.90751 V/mu_s
** Phase margin: 60.1606°
** CMRR: 141 dB
** VoutMax: 4.25 V
** VoutMin: 1.60001 V
** VcmMax: 5.11001 V
** VcmMin: 1.42001 V


** Expected Currents: 
** NormalTransistorPmos: -2.24369e+07 muA
** NormalTransistorPmos: -4.02299e+07 muA
** NormalTransistorPmos: -2.38002e+08 muA
** NormalTransistorPmos: -2.24389e+07 muA
** NormalTransistorPmos: -3.69579e+07 muA
** NormalTransistorPmos: -2.24389e+07 muA
** NormalTransistorPmos: -3.69579e+07 muA
** DiodeTransistorNmos: 2.24381e+07 muA
** NormalTransistorNmos: 2.24381e+07 muA
** NormalTransistorNmos: 2.24381e+07 muA
** NormalTransistorNmos: 2.90351e+07 muA
** DiodeTransistorNmos: 2.90341e+07 muA
** NormalTransistorNmos: 1.45181e+07 muA
** NormalTransistorNmos: 1.45181e+07 muA
** NormalTransistorNmos: 1.87331e+09 muA
** DiodeTransistorNmos: 1.87331e+09 muA
** NormalTransistorPmos: -1.8733e+09 muA
** DiodeTransistorNmos: 2.24361e+07 muA
** NormalTransistorNmos: 2.24351e+07 muA
** DiodeTransistorNmos: 4.02291e+07 muA
** NormalTransistorNmos: 4.02301e+07 muA
** DiodeTransistorNmos: 2.38003e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.18001  V
** outInputVoltageBiasXXnXX2: 2.01001  V
** outSourceVoltageBiasXXnXX1: 0.590001  V
** outSourceVoltageBiasXXnXX2: 1.00501  V
** outSourceVoltageBiasXXpXX1: 4.13601  V
** outVoltageBiasXXnXX3: 0.983001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.407001  V
** out1: 0.612001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.85501  V
** inner: 0.589001  V
** inner: 1.00601  V


.END