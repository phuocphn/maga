** Name: two_stage_single_output_op_amp_96_12

.MACRO two_stage_single_output_op_amp_96_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=98e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=163e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=141e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=237e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mTelescopicFirstStageLoad7 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=63e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=74e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=74e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=98e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=163e-6
mTelescopicFirstStageLoad12 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=63e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=119e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=233e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=282e-6
mTelescopicFirstStageLoad16 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=37e-6
mTelescopicFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=32e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=32e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=560e-6
mMainBias20 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=482e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=489e-6
mTelescopicFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=37e-6
mMainBias23 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=463e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.2001e-12
.EOM two_stage_single_output_op_amp_96_12

** Expected Performance Values: 
** Gain: 200 dB
** Power consumption: 4.97501 mW
** Area: 10300 (mu_m)^2
** Transit frequency: 3.49501 MHz
** Transit frequency with error factor: 3.49452 MHz
** Slew rate: 9.599 V/mu_s
** Phase margin: 60.1606°
** CMRR: 130 dB
** VoutMax: 4.64001 V
** VoutMin: 0.700001 V
** VcmMax: 4.72001 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 9.19981e+07 muA
** NormalTransistorNmos: 1.78401e+08 muA
** NormalTransistorPmos: -1.86654e+08 muA
** NormalTransistorPmos: -1.77263e+08 muA
** NormalTransistorNmos: 2.01361e+07 muA
** NormalTransistorNmos: 2.01341e+07 muA
** NormalTransistorPmos: -2.01369e+07 muA
** NormalTransistorPmos: -2.01359e+07 muA
** NormalTransistorPmos: -2.01349e+07 muA
** NormalTransistorPmos: -2.01359e+07 muA
** NormalTransistorNmos: 2.17533e+08 muA
** NormalTransistorNmos: 2.01351e+07 muA
** NormalTransistorNmos: 2.01351e+07 muA
** NormalTransistorNmos: 3.10455e+08 muA
** DiodeTransistorNmos: 3.10455e+08 muA
** NormalTransistorPmos: -3.10454e+08 muA
** NormalTransistorPmos: -3.10455e+08 muA
** DiodeTransistorNmos: 1.86655e+08 muA
** NormalTransistorNmos: 1.86655e+08 muA
** DiodeTransistorNmos: 1.77264e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.19989e+07 muA
** DiodeTransistorPmos: -1.784e+08 muA


** Expected Voltages: 
** ibias: 0.570001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11001  V
** out: 2.5  V
** outFirstStage: 4.25901  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 4.18201  V
** outVoltageBiasXXpXX1: 3.69501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 3.90301  V
** innerTransistorStack1Load2: 4.43301  V
** innerTransistorStack2Load2: 4.43301  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.44701  V
** inner: 0.555001  V


.END