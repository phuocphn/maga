** Name: one_stage_single_output_op_amp80

.MACRO one_stage_single_output_op_amp80 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=67e-6
mFoldedCascodeFirstStageStageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=64e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=14e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=239e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=65e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=65e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=44e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=44e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=64e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=67e-6
mFoldedCascodeFirstStageLoad13 out outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=239e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=130e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=185e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=185e-6
mFoldedCascodeFirstStageLoad17 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=130e-6
mMainBias18 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=130e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp80

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 2.74001 mW
** Area: 4962 (mu_m)^2
** Transit frequency: 4.41601 MHz
** Transit frequency with error factor: 4.41564 MHz
** Slew rate: 6.22593 V/mu_s
** Phase margin: 88.8085°
** CMRR: 142 dB
** VoutMax: 3.97001 V
** VoutMin: 0.310001 V
** VcmMax: 5.17001 V
** VcmMin: 1.83001 V


** Expected Currents: 
** NormalTransistorPmos: -1.30945e+08 muA
** NormalTransistorPmos: -2.19789e+07 muA
** NormalTransistorPmos: -1.25042e+08 muA
** NormalTransistorPmos: -1.87562e+08 muA
** NormalTransistorPmos: -1.25046e+08 muA
** NormalTransistorPmos: -1.87566e+08 muA
** NormalTransistorNmos: 1.25045e+08 muA
** NormalTransistorNmos: 1.25046e+08 muA
** NormalTransistorNmos: 1.25047e+08 muA
** NormalTransistorNmos: 1.25046e+08 muA
** NormalTransistorNmos: 1.25042e+08 muA
** DiodeTransistorNmos: 1.25041e+08 muA
** NormalTransistorNmos: 6.25211e+07 muA
** NormalTransistorNmos: 6.25211e+07 muA
** DiodeTransistorNmos: 1.30946e+08 muA
** NormalTransistorNmos: 1.30945e+08 muA
** DiodeTransistorNmos: 2.19781e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.43501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outInputVoltageBiasXXnXX1: 1.61001  V
** outSourceVoltageBiasXXnXX1: 0.805001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.912001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 4.23001  V
** sourceGCC2: 4.23001  V
** sourceTransconductance: 1.87001  V
** inner: 0.801001  V


.END