** Name: two_stage_single_output_op_amp_197_9

.MACRO two_stage_single_output_op_amp_197_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=4e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=7e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=7e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=99e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=32e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=81e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=12e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=23e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=15e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=46e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=99e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=4e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=15e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=60e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=60e-6
mSimpleFirstStageLoad19 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=6e-6 W=600e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=31e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=171e-6
mSimpleFirstStageLoad22 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=600e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=72e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_197_9

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 5.38001 mW
** Area: 11408 (mu_m)^2
** Transit frequency: 4.29601 MHz
** Transit frequency with error factor: 4.29345 MHz
** Slew rate: 4.04866 V/mu_s
** Phase margin: 63.0254°
** CMRR: 109 dB
** VoutMax: 4.25 V
** VoutMin: 1.84001 V
** VcmMax: 4.71001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorPmos: -6.06269e+07 muA
** NormalTransistorPmos: -2.62949e+07 muA
** DiodeTransistorNmos: 4.09501e+07 muA
** DiodeTransistorNmos: 4.09511e+07 muA
** NormalTransistorNmos: 4.09501e+07 muA
** NormalTransistorNmos: 4.09511e+07 muA
** NormalTransistorPmos: -5.04749e+07 muA
** NormalTransistorPmos: -5.04759e+07 muA
** NormalTransistorPmos: -5.04749e+07 muA
** NormalTransistorPmos: -5.04759e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90461e+07 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 8.68116e+08 muA
** DiodeTransistorNmos: 8.68115e+08 muA
** NormalTransistorPmos: -8.68115e+08 muA
** DiodeTransistorNmos: 6.06261e+07 muA
** NormalTransistorNmos: 6.06251e+07 muA
** DiodeTransistorNmos: 2.62941e+07 muA
** DiodeTransistorNmos: 2.62931e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.62601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 2.24401  V
** outSourceVoltageBiasXXnXX1: 1.12201  V
** outSourceVoltageBiasXXnXX2: 0.666001  V
** outSourceVoltageBiasXXpXX1: 3.90501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.10401  V
** innerStageBias: 1.03601  V
** innerTransistorStack1Load2: 3.86901  V
** innerTransistorStack2Load1: 1.10401  V
** innerTransistorStack2Load2: 3.86901  V
** out1: 2.20701  V
** sourceTransconductance: 1.94501  V
** inner: 1.12101  V


.END