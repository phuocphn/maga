** Name: two_stage_single_output_op_amp_87_2

.MACRO two_stage_single_output_op_amp_87_2 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=199e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=94e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=15e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=199e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=213e-6
mMainBias8 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=128e-6
mSecondStage1Transconductor9 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=428e-6
mTelescopicFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=57e-6
mTelescopicFirstStageLoad11 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=4e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=76e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=76e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mSecondStage1StageBias15 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mTelescopicFirstStageLoad16 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=4e-6
mMainBias17 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=311e-6
mTelescopicFirstStageStageBias18 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=594e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.1001e-12
.EOM two_stage_single_output_op_amp_87_2

** Expected Performance Values: 
** Gain: 135 dB
** Power consumption: 5.30801 mW
** Area: 6223 (mu_m)^2
** Transit frequency: 5.71901 MHz
** Transit frequency with error factor: 5.71917 MHz
** Slew rate: 11.5432 V/mu_s
** Phase margin: 60.1606°
** CMRR: 124 dB
** VoutMax: 4.81001 V
** VoutMin: 0.300001 V
** VcmMax: 4.04001 V
** VcmMin: 1.89001 V


** Expected Currents: 
** NormalTransistorNmos: 2.92007e+08 muA
** NormalTransistorPmos: -2.10198e+08 muA
** NormalTransistorPmos: -2.30869e+07 muA
** NormalTransistorPmos: -5.43689e+07 muA
** NormalTransistorPmos: -5.43689e+07 muA
** DiodeTransistorNmos: 5.43681e+07 muA
** NormalTransistorNmos: 5.43681e+07 muA
** NormalTransistorNmos: 5.43681e+07 muA
** NormalTransistorPmos: -4.00743e+08 muA
** NormalTransistorPmos: -5.43679e+07 muA
** NormalTransistorPmos: -5.43679e+07 muA
** NormalTransistorNmos: 4.07609e+08 muA
** NormalTransistorNmos: 4.07608e+08 muA
** NormalTransistorPmos: -4.07608e+08 muA
** DiodeTransistorNmos: 2.10199e+08 muA
** DiodeTransistorNmos: 2.30861e+07 muA
** DiodeTransistorPmos: -2.92006e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXpXX1: 0.623001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.636001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.26401  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 2.93901  V
** sourceGCC2: 2.93901  V
** innerTransconductance: 0.150001  V


.END