** Name: two_stage_single_output_op_amp_190_10

.MACRO two_stage_single_output_op_amp_190_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=268e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=6e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=113e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=121e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=268e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=113e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=6e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=554e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=46e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=121e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=40e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=599e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=599e-6
mSimpleFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=359e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=496e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=359e-6
mMainBias22 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.8001e-12
.EOM two_stage_single_output_op_amp_190_10

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 14.9991 mW
** Area: 14310 (mu_m)^2
** Transit frequency: 8.76901 MHz
** Transit frequency with error factor: 8.76436 MHz
** Slew rate: 8.26487 V/mu_s
** Phase margin: 60.1606°
** CMRR: 116 dB
** VoutMax: 4.25 V
** VoutMin: 0.340001 V
** VcmMax: 4.69001 V
** VcmMin: 1.45001 V


** Expected Currents: 
** NormalTransistorNmos: 9.95231e+07 muA
** NormalTransistorNmos: 9.80301e+06 muA
** NormalTransistorPmos: -6.12199e+06 muA
** NormalTransistorNmos: 6.89456e+08 muA
** NormalTransistorNmos: 6.89456e+08 muA
** DiodeTransistorNmos: 6.89456e+08 muA
** NormalTransistorPmos: -7.4707e+08 muA
** NormalTransistorPmos: -7.47069e+08 muA
** NormalTransistorPmos: -7.4707e+08 muA
** NormalTransistorPmos: -7.47069e+08 muA
** NormalTransistorNmos: 1.1523e+08 muA
** DiodeTransistorNmos: 1.15229e+08 muA
** NormalTransistorNmos: 5.76151e+07 muA
** NormalTransistorNmos: 5.76151e+07 muA
** NormalTransistorNmos: 1.38032e+09 muA
** NormalTransistorPmos: -1.38031e+09 muA
** NormalTransistorPmos: -1.38031e+09 muA
** DiodeTransistorNmos: 6.12101e+06 muA
** NormalTransistorNmos: 6.12001e+06 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.95239e+07 muA
** DiodeTransistorPmos: -9.80199e+06 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.04301  V
** outInputVoltageBiasXXnXX1: 1.30001  V
** outSourceVoltageBiasXXnXX1: 0.650001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.06401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.59001  V
** innerTransistorStack2Load1: 0.958001  V
** innerTransistorStack2Load2: 4.59001  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.60701  V
** inner: 0.649001  V


.END