** Name: two_stage_single_output_op_amp_94_7

.MACRO two_stage_single_output_op_amp_94_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=83e-6
mTelescopicFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=31e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=8e-6
mTelescopicFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=9e-6 W=29e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=29e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=29e-6
mMainBias9 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=33e-6
mSecondStage1StageBias10 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=9e-6 W=29e-6
mMainBias12 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mTelescopicFirstStageStageBias13 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=67e-6
mTelescopicFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=31e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=516e-6
mTelescopicFirstStageLoad16 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=25e-6
mMainBias17 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=77e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_94_7

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 4.45101 mW
** Area: 5530 (mu_m)^2
** Transit frequency: 2.88501 MHz
** Transit frequency with error factor: 2.88453 MHz
** Slew rate: 18.183 V/mu_s
** Phase margin: 64.1713°
** CMRR: 134 dB
** VoutMax: 4.5 V
** VoutMin: 0.170001 V
** VcmMax: 4.22001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorNmos: 7.37401e+06 muA
** NormalTransistorNmos: 4.05621e+07 muA
** NormalTransistorPmos: -6.98259e+07 muA
** NormalTransistorNmos: 6.13901e+06 muA
** NormalTransistorNmos: 6.13801e+06 muA
** DiodeTransistorPmos: -6.13999e+06 muA
** NormalTransistorPmos: -6.13899e+06 muA
** NormalTransistorPmos: -6.13999e+06 muA
** NormalTransistorNmos: 8.21001e+07 muA
** NormalTransistorNmos: 6.13801e+06 muA
** NormalTransistorNmos: 6.13801e+06 muA
** NormalTransistorNmos: 7.50076e+08 muA
** NormalTransistorPmos: -7.50075e+08 muA
** DiodeTransistorNmos: 6.98251e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.375e+06 muA
** DiodeTransistorPmos: -4.05629e+07 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.37601  V
** out: 2.5  V
** outFirstStage: 3.94001  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 3.98401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 4.20101  V
** out1: 4.22501  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END