** Name: two_stage_single_output_op_amp_79_10

.MACRO two_stage_single_output_op_amp_79_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=48e-6
mMainBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageStageBias5 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=79e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=171e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=9e-6 W=207e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=171e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=277e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=96e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=92e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=482e-6
mMainBias20 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=48e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=448e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=92e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_79_10

** Expected Performance Values: 
** Gain: 141 dB
** Power consumption: 4.17501 mW
** Area: 10939 (mu_m)^2
** Transit frequency: 5.29401 MHz
** Transit frequency with error factor: 5.2938 MHz
** Slew rate: 4.0782 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.59001 V
** VoutMin: 0.170001 V
** VcmMax: 5.01001 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorNmos: 1.62454e+08 muA
** NormalTransistorNmos: 5.57561e+07 muA
** NormalTransistorPmos: -1.33817e+08 muA
** NormalTransistorPmos: -3.73639e+07 muA
** NormalTransistorPmos: -6.02209e+07 muA
** NormalTransistorPmos: -3.73639e+07 muA
** NormalTransistorPmos: -6.02209e+07 muA
** NormalTransistorNmos: 3.73631e+07 muA
** NormalTransistorNmos: 3.73621e+07 muA
** NormalTransistorNmos: 3.73631e+07 muA
** NormalTransistorNmos: 3.73621e+07 muA
** NormalTransistorNmos: 4.57111e+07 muA
** NormalTransistorNmos: 4.57101e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 3.52437e+08 muA
** NormalTransistorPmos: -3.52436e+08 muA
** NormalTransistorPmos: -3.52437e+08 muA
** DiodeTransistorNmos: 1.33818e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.62453e+08 muA
** DiodeTransistorPmos: -5.57569e+07 muA


** Expected Voltages: 
** ibias: 0.571001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.948001  V
** out: 2.5  V
** outFirstStage: 4.23301  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.04301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.390001  V
** innerTransistorStack1Load2: 0.390001  V
** innerTransistorStack2Load2: 0.391001  V
** out1: 0.596001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.45901  V


.END