** Name: two_stage_single_output_op_amp_138_6

.MACRO two_stage_single_output_op_amp_138_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=21e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=4e-6 W=10e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=10e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=120e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=12e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=93e-6
mSimpleFirstStageLoad8 FirstStageYinnerOutputLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=73e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=100e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=100e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=87e-6
mSecondStage1Transconductor12 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=208e-6
mSimpleFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=73e-6
mMainBias14 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=43e-6
mSimpleFirstStageTransconductor15 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=125e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=10e-6
mSimpleFirstStageStageBias17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=7e-6 W=600e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=12e-6
mMainBias19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=282e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=124e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=93e-6
mSimpleFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=10e-6
mSimpleFirstStageTransconductor23 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=125e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.70001e-12
.EOM two_stage_single_output_op_amp_138_6

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 1.71201 mW
** Area: 14775 (mu_m)^2
** Transit frequency: 2.58801 MHz
** Transit frequency with error factor: 2.58529 MHz
** Slew rate: 5.196 V/mu_s
** Phase margin: 60.1606°
** CMRR: 86 dB
** VoutMax: 3.17001 V
** VoutMin: 0.340001 V
** VcmMax: 3.94001 V
** VcmMin: -0.159999 V


** Expected Currents: 
** NormalTransistorNmos: 2.14101e+07 muA
** NormalTransistorPmos: -2.33519e+07 muA
** NormalTransistorPmos: -1.04569e+07 muA
** DiodeTransistorPmos: -2.53829e+07 muA
** NormalTransistorPmos: -2.53829e+07 muA
** NormalTransistorPmos: -2.53829e+07 muA
** DiodeTransistorPmos: -2.53829e+07 muA
** NormalTransistorNmos: 5.07261e+07 muA
** NormalTransistorNmos: 5.07251e+07 muA
** NormalTransistorNmos: 5.07261e+07 muA
** NormalTransistorNmos: 5.07251e+07 muA
** NormalTransistorPmos: -5.06869e+07 muA
** NormalTransistorPmos: -2.53439e+07 muA
** NormalTransistorPmos: -2.53439e+07 muA
** NormalTransistorNmos: 1.65703e+08 muA
** NormalTransistorNmos: 1.65704e+08 muA
** NormalTransistorPmos: -1.65702e+08 muA
** DiodeTransistorPmos: -1.65703e+08 muA
** DiodeTransistorNmos: 2.33511e+07 muA
** DiodeTransistorNmos: 1.04561e+07 muA
** DiodeTransistorPmos: -2.14109e+07 muA
** NormalTransistorPmos: -2.14119e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.804001  V
** inputVoltageBiasXXnXX2: 0.623001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.60401  V
** outSourceVoltageBiasXXpXX1: 3.80201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.218001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.218001  V
** sourceTransconductance: 3.38201  V
** innerTransconductance: 0.205001  V
** inner: 3.79701  V


.END