** Name: symmetrical_op_amp185

.MACRO symmetrical_op_amp185 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=2e-6 W=35e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias5 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=106e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=34e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=40e-6
mSecondStage1StageBias10 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=58e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=40e-6
mMainBias12 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=207e-6
mSymmetricalFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=20e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=20e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=44e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=44e-6
mSymmetricalFirstStageLoad17 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=63e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=141e-6
mSecondStage1Transconductor19 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=141e-6
mSymmetricalFirstStageLoad20 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=63e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp185

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 1.37201 mW
** Area: 3040 (mu_m)^2
** Transit frequency: 5.91501 MHz
** Transit frequency with error factor: 5.91479 MHz
** Slew rate: 5.6866 V/mu_s
** Phase margin: 79.6412°
** CMRR: 145 dB
** negPSRR: 124 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 0.910001 V
** VcmMax: 4.81001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 9.95591e+07 muA
** NormalTransistorPmos: -2.53969e+07 muA
** NormalTransistorPmos: -2.53979e+07 muA
** NormalTransistorPmos: -2.53969e+07 muA
** NormalTransistorPmos: -2.53979e+07 muA
** NormalTransistorNmos: 5.07911e+07 muA
** NormalTransistorNmos: 5.07901e+07 muA
** NormalTransistorNmos: 2.53961e+07 muA
** NormalTransistorNmos: 2.53961e+07 muA
** NormalTransistorNmos: 5.69931e+07 muA
** NormalTransistorNmos: 5.69921e+07 muA
** NormalTransistorPmos: -5.69939e+07 muA
** NormalTransistorPmos: -5.69929e+07 muA
** DiodeTransistorNmos: 5.69911e+07 muA
** DiodeTransistorNmos: 5.69901e+07 muA
** NormalTransistorPmos: -5.69919e+07 muA
** NormalTransistorPmos: -5.69929e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -9.95599e+07 muA


** Expected Voltages: 
** ibias: 1.17701  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 0.754001  V
** inSourceTransconductanceComplementarySecondStage: 3.83701  V
** innerComplementarySecondStage: 1.35501  V
** out: 2.5  V
** out1FirstStage: 3.83701  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.505001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.797001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END