** Name: two_stage_single_output_op_amp_143_12

.MACRO two_stage_single_output_op_amp_143_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=27e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=19e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=9e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=300e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=5e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=300e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=27e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=217e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
mMainBias11 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=29e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=300e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=15e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=300e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=462e-6
mSimpleFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=53e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=484e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=53e-6
mMainBias20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=13e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.7001e-12
.EOM two_stage_single_output_op_amp_143_12

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 9.98001 mW
** Area: 14984 (mu_m)^2
** Transit frequency: 6.45401 MHz
** Transit frequency with error factor: 6.44202 MHz
** Slew rate: 6.08273 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 1.20001 V
** VcmMax: 4.69001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorNmos: 2.43681e+08 muA
** NormalTransistorNmos: 1.52841e+07 muA
** NormalTransistorPmos: -4.04359e+07 muA
** NormalTransistorNmos: 1.07545e+08 muA
** NormalTransistorNmos: 1.07545e+08 muA
** DiodeTransistorNmos: 1.07545e+08 muA
** NormalTransistorPmos: -1.64683e+08 muA
** NormalTransistorPmos: -1.64683e+08 muA
** NormalTransistorNmos: 1.14278e+08 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 1.35721e+09 muA
** DiodeTransistorNmos: 1.35721e+09 muA
** NormalTransistorPmos: -1.3572e+09 muA
** NormalTransistorPmos: -1.35721e+09 muA
** DiodeTransistorNmos: 4.04351e+07 muA
** NormalTransistorNmos: 4.04341e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.4368e+08 muA
** DiodeTransistorPmos: -1.52849e+07 muA


** Expected Voltages: 
** ibias: 0.613001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.71701  V
** out: 2.5  V
** outFirstStage: 4.04001  V
** outInputVoltageBiasXXnXX1: 1.60801  V
** outSourceVoltageBiasXXnXX1: 0.804001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 1.05901  V
** out1: 2.11801  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.60401  V
** inner: 0.802001  V


.END