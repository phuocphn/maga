** Name: two_stage_single_output_op_amp_148_10

.MACRO two_stage_single_output_op_amp_148_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=41e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=2e-6 W=22e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=139e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=341e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=9e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=2e-6 W=22e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=63e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=448e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=41e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=9e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mMainBias13 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=427e-6
mSimpleFirstStageLoad14 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=342e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=567e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=567e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=565e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=351e-6
mSimpleFirstStageLoad19 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=342e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.10001e-12
.EOM two_stage_single_output_op_amp_148_10

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 11.0251 mW
** Area: 11651 (mu_m)^2
** Transit frequency: 3.44501 MHz
** Transit frequency with error factor: 3.44049 MHz
** Slew rate: 6.64888 V/mu_s
** Phase margin: 60.1606°
** CMRR: 116 dB
** VoutMax: 4.28001 V
** VoutMin: 0.160001 V
** VcmMax: 4.67001 V
** VcmMin: 0.880001 V


** Expected Currents: 
** NormalTransistorNmos: 4.65575e+08 muA
** NormalTransistorNmos: 3.25611e+08 muA
** DiodeTransistorNmos: 5.07582e+08 muA
** DiodeTransistorNmos: 5.07583e+08 muA
** NormalTransistorNmos: 5.07582e+08 muA
** NormalTransistorNmos: 5.07583e+08 muA
** NormalTransistorPmos: -5.3154e+08 muA
** NormalTransistorPmos: -5.31541e+08 muA
** NormalTransistorPmos: -5.3154e+08 muA
** NormalTransistorPmos: -5.31541e+08 muA
** NormalTransistorNmos: 4.79181e+07 muA
** NormalTransistorNmos: 2.39591e+07 muA
** NormalTransistorNmos: 2.39591e+07 muA
** NormalTransistorNmos: 3.40747e+08 muA
** NormalTransistorPmos: -3.40746e+08 muA
** NormalTransistorPmos: -3.40747e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.65574e+08 muA
** DiodeTransistorPmos: -3.2561e+08 muA


** Expected Voltages: 
** ibias: 0.570001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.11701  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.20601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerTransistorStack1Load1: 1.14701  V
** innerTransistorStack1Load2: 4.75901  V
** innerTransistorStack2Load1: 1.14701  V
** innerTransistorStack2Load2: 4.75901  V
** sourceTransconductance: 1.78701  V
** innerTransconductance: 4.65201  V


.END