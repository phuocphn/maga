** Name: two_stage_single_output_op_amp_60_1

.MACRO two_stage_single_output_op_amp_60_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=14e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=93e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=61e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=128e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=22e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=65e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=65e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=332e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=22e-6
mMainBias12 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=62e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=93e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=53e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=53e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=128e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=61e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=566e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=43e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_60_1

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 4.95001 mW
** Area: 8327 (mu_m)^2
** Transit frequency: 4.04401 MHz
** Transit frequency with error factor: 4.04426 MHz
** Slew rate: 4.54435 V/mu_s
** Phase margin: 71.0468°
** CMRR: 144 dB
** VoutMax: 4.58001 V
** VoutMin: 0.530001 V
** VcmMax: 3.22001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.00001e+07 muA
** NormalTransistorNmos: 2.98191e+07 muA
** NormalTransistorNmos: 2.05231e+07 muA
** NormalTransistorNmos: 3.09511e+07 muA
** NormalTransistorNmos: 2.05231e+07 muA
** NormalTransistorNmos: 3.09511e+07 muA
** NormalTransistorPmos: -2.05239e+07 muA
** NormalTransistorPmos: -2.05239e+07 muA
** DiodeTransistorPmos: -2.05239e+07 muA
** NormalTransistorPmos: -2.08589e+07 muA
** DiodeTransistorPmos: -2.08599e+07 muA
** NormalTransistorPmos: -1.04289e+07 muA
** NormalTransistorPmos: -1.04289e+07 muA
** NormalTransistorNmos: 8.78327e+08 muA
** NormalTransistorPmos: -8.78326e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.00009e+07 muA
** NormalTransistorPmos: -1.00019e+07 muA
** DiodeTransistorPmos: -2.98199e+07 muA


** Expected Voltages: 
** ibias: 1.14301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.938001  V
** outInputVoltageBiasXXpXX1: 3.40201  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.20101  V
** outVoltageBiasXXpXX2: 4.01801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.27901  V
** out1: 3.55101  V
** sourceGCC1: 0.527001  V
** sourceGCC2: 0.527001  V
** sourceTransconductance: 3.24501  V
** inner: 4.20001  V


.END