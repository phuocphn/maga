** Name: two_stage_single_output_op_amp_169_4

.MACRO two_stage_single_output_op_amp_169_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=88e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=553e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=528e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=74e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=39e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSimpleFirstStageLoad7 FirstStageYinnerOutputLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=505e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=487e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=487e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=297e-6
mSecondStage1Transconductor11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=286e-6
mSimpleFirstStageLoad12 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=505e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=361e-6
mSimpleFirstStageStageBias14 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=25e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=74e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=100e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=139e-6
mSecondStage1StageBias18 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=600e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=528e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=361e-6
mMainBias21 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=168e-6
mMainBias22 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=266e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.30001e-12
.EOM two_stage_single_output_op_amp_169_4

** Expected Performance Values: 
** Gain: 152 dB
** Power consumption: 10.7431 mW
** Area: 14636 (mu_m)^2
** Transit frequency: 5.45101 MHz
** Transit frequency with error factor: 5.44712 MHz
** Slew rate: 5.26946 V/mu_s
** Phase margin: 60.1606°
** CMRR: 127 dB
** VoutMax: 3.73001 V
** VoutMin: 0.300001 V
** VcmMax: 3.01001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorPmos: -3.42101e+08 muA
** NormalTransistorPmos: -5.4166e+08 muA
** DiodeTransistorPmos: -4.55463e+08 muA
** DiodeTransistorPmos: -4.55464e+08 muA
** NormalTransistorPmos: -4.55463e+08 muA
** NormalTransistorPmos: -4.55464e+08 muA
** NormalTransistorNmos: 4.80919e+08 muA
** NormalTransistorNmos: 4.80918e+08 muA
** NormalTransistorNmos: 4.80919e+08 muA
** NormalTransistorNmos: 4.80918e+08 muA
** NormalTransistorPmos: -5.09089e+07 muA
** NormalTransistorPmos: -5.09079e+07 muA
** NormalTransistorPmos: -2.54549e+07 muA
** NormalTransistorPmos: -2.54549e+07 muA
** NormalTransistorNmos: 2.83049e+08 muA
** NormalTransistorNmos: 2.83048e+08 muA
** NormalTransistorPmos: -2.83048e+08 muA
** NormalTransistorPmos: -2.83047e+08 muA
** DiodeTransistorNmos: 3.42102e+08 muA
** DiodeTransistorNmos: 5.41661e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.22701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.96101  V
** outVoltageBiasXXnXX1: 0.708001  V
** outVoltageBiasXXnXX2: 0.557001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.06301  V
** innerSourceLoad1: 3.84701  V
** innerStageBias: 4.02901  V
** innerTransistorStack1Load2: 0.153001  V
** innerTransistorStack2Load1: 3.84601  V
** innerTransistorStack2Load2: 0.153001  V
** sourceTransconductance: 3.21801  V
** innerStageBias: 4.02001  V
** innerTransconductance: 0.150001  V


.END