** Name: one_stage_single_output_op_amp109

.MACRO one_stage_single_output_op_amp109 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=41e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=41e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=26e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=18e-6
mMainBias5 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=10e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=41e-6
mTelescopicFirstStageLoad8 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=41e-6
mMainBias9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=42e-6
mTelescopicFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=56e-6
mTelescopicFirstStageLoad11 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=38e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=154e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=154e-6
mTelescopicFirstStageLoad14 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=38e-6
mMainBias15 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=567e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp109

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 0.762001 mW
** Area: 3758 (mu_m)^2
** Transit frequency: 2.71501 MHz
** Transit frequency with error factor: 2.71533 MHz
** Slew rate: 5.69573 V/mu_s
** Phase margin: 85.9437°
** CMRR: 140 dB
** VoutMax: 3.07001 V
** VoutMin: 0.720001 V
** VcmMax: 3 V
** VcmMin: 1.06001 V


** Expected Currents: 
** NormalTransistorNmos: 2.92411e+07 muA
** NormalTransistorPmos: -1.83259e+07 muA
** NormalTransistorPmos: -4.23979e+07 muA
** NormalTransistorPmos: -4.23979e+07 muA
** DiodeTransistorNmos: 4.23971e+07 muA
** NormalTransistorNmos: 4.23961e+07 muA
** NormalTransistorNmos: 4.23971e+07 muA
** DiodeTransistorNmos: 4.23961e+07 muA
** NormalTransistorPmos: -1.14034e+08 muA
** NormalTransistorPmos: -1.14033e+08 muA
** NormalTransistorPmos: -4.23969e+07 muA
** NormalTransistorPmos: -4.23969e+07 muA
** DiodeTransistorNmos: 1.83251e+07 muA
** DiodeTransistorPmos: -2.92419e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.14701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX2: 3.96101  V
** outVoltageBiasXXnXX0: 0.662001  V
** outVoltageBiasXXpXX1: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.31101  V
** innerSourceLoad2: 0.561001  V
** innerStageBias: 3.86101  V
** innerTransistorStack1Load2: 0.560001  V
** out1: 1.12201  V
** sourceGCC1: 2.99901  V
** sourceGCC2: 2.99901  V


.END