** Name: two_stage_single_output_op_amp_68_3

.MACRO two_stage_single_output_op_amp_68_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=32e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=33e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=33e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=17e-6
mMainBias6 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=6e-6 W=9e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=144e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=11e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=40e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=88e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=88e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=10e-6 W=223e-6
mFoldedCascodeFirstStageLoad13 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=40e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias15 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=51e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=33e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=112e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=112e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=144e-6
mSecondStage1StageBias20 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=388e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=17e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=6e-6 W=316e-6
mFoldedCascodeFirstStageLoad23 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=33e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_68_3

** Expected Performance Values: 
** Gain: 131 dB
** Power consumption: 2.81101 mW
** Area: 12782 (mu_m)^2
** Transit frequency: 3.18101 MHz
** Transit frequency with error factor: 3.18078 MHz
** Slew rate: 3.50834 V/mu_s
** Phase margin: 61.3065°
** CMRR: 145 dB
** VoutMax: 3.07001 V
** VoutMin: 0.510001 V
** VcmMax: 3.34001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.91101e+06 muA
** NormalTransistorNmos: 1.41081e+07 muA
** NormalTransistorNmos: 1.58641e+07 muA
** NormalTransistorNmos: 2.40241e+07 muA
** NormalTransistorNmos: 1.58641e+07 muA
** NormalTransistorNmos: 2.40241e+07 muA
** DiodeTransistorPmos: -1.58649e+07 muA
** NormalTransistorPmos: -1.58659e+07 muA
** NormalTransistorPmos: -1.58649e+07 muA
** DiodeTransistorPmos: -1.58659e+07 muA
** NormalTransistorPmos: -1.63229e+07 muA
** DiodeTransistorPmos: -1.63239e+07 muA
** NormalTransistorPmos: -8.16099e+06 muA
** NormalTransistorPmos: -8.16099e+06 muA
** NormalTransistorNmos: 4.88038e+08 muA
** NormalTransistorPmos: -4.88037e+08 muA
** NormalTransistorPmos: -4.88038e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.91199e+06 muA
** NormalTransistorPmos: -1.91299e+06 muA
** DiodeTransistorPmos: -1.41089e+07 muA
** DiodeTransistorPmos: -1.41099e+07 muA


** Expected Voltages: 
** ibias: 1.12101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.916001  V
** outInputVoltageBiasXXpXX1: 3.51601  V
** outInputVoltageBiasXXpXX2: 2.49001  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outSourceVoltageBiasXXpXX1: 4.25801  V
** outSourceVoltageBiasXXpXX2: 3.78301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.27201  V
** innerTransistorStack2Load2: 4.27201  V
** out1: 3.54401  V
** sourceGCC1: 0.534001  V
** sourceGCC2: 0.534001  V
** sourceTransconductance: 3.24401  V
** innerStageBias: 3.77101  V
** inner: 4.25701  V


.END