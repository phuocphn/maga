** Name: two_stage_single_output_op_amp_74_9

.MACRO two_stage_single_output_op_amp_74_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=31e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=28e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=8e-6 W=8e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=181e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=41e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=23e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=31e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=12e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=12e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=28e-6
mMainBias13 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=8e-6 W=181e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=3e-6 W=10e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=160e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=58e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=58e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=213e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=160e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=99e-6
mMainBias22 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=105e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_74_9

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 6.13101 mW
** Area: 6934 (mu_m)^2
** Transit frequency: 2.58201 MHz
** Transit frequency with error factor: 2.58207 MHz
** Slew rate: 3.56892 V/mu_s
** Phase margin: 66.4632°
** CMRR: 139 dB
** VoutMax: 4.25 V
** VoutMin: 1.89001 V
** VcmMax: 5.09001 V
** VcmMin: 1.45001 V


** Expected Currents: 
** NormalTransistorPmos: -4.32549e+07 muA
** NormalTransistorPmos: -4.64199e+07 muA
** NormalTransistorPmos: -1.62449e+07 muA
** NormalTransistorPmos: -2.56409e+07 muA
** NormalTransistorPmos: -1.62449e+07 muA
** NormalTransistorPmos: -2.56409e+07 muA
** NormalTransistorNmos: 1.62441e+07 muA
** NormalTransistorNmos: 1.62441e+07 muA
** DiodeTransistorNmos: 1.62441e+07 muA
** NormalTransistorNmos: 1.87891e+07 muA
** DiodeTransistorNmos: 1.87881e+07 muA
** NormalTransistorNmos: 9.39501e+06 muA
** NormalTransistorNmos: 9.39501e+06 muA
** NormalTransistorNmos: 1.06528e+09 muA
** DiodeTransistorNmos: 1.06528e+09 muA
** NormalTransistorPmos: -1.06527e+09 muA
** DiodeTransistorNmos: 4.32541e+07 muA
** NormalTransistorNmos: 4.32551e+07 muA
** DiodeTransistorNmos: 4.64191e+07 muA
** NormalTransistorNmos: 4.64181e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.19401  V
** outInputVoltageBiasXXnXX2: 2.29601  V
** outSourceVoltageBiasXXnXX1: 0.597001  V
** outSourceVoltageBiasXXnXX2: 1.14801  V
** outSourceVoltageBiasXXpXX1: 4.12301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.581001  V
** out1: 1.22501  V
** sourceGCC1: 4.03901  V
** sourceGCC2: 4.03901  V
** sourceTransconductance: 1.84001  V
** inner: 0.598001  V
** inner: 1.14701  V


.END