** Name: two_stage_single_output_op_amp_39_9

.MACRO two_stage_single_output_op_amp_39_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=17e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=474e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=27e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=5e-6 W=27e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=9e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=59e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=15e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=47e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=16e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=474e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=15e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=27e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=456e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=27e-6
mMainBias18 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=30e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_39_9

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 3.50301 mW
** Area: 8091 (mu_m)^2
** Transit frequency: 4.11401 MHz
** Transit frequency with error factor: 4.11153 MHz
** Slew rate: 3.87762 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** negPSRR: 101 dB
** posPSRR: 94 dB
** VoutMax: 4.25 V
** VoutMin: 0.840001 V
** VcmMax: 3.62001 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorNmos: 5.18601e+06 muA
** NormalTransistorPmos: -1.75809e+07 muA
** DiodeTransistorPmos: -9.52499e+06 muA
** NormalTransistorPmos: -9.52599e+06 muA
** NormalTransistorPmos: -9.52499e+06 muA
** DiodeTransistorPmos: -9.52599e+06 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90461e+07 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 6.48734e+08 muA
** DiodeTransistorNmos: 6.48733e+08 muA
** NormalTransistorPmos: -6.48733e+08 muA
** DiodeTransistorNmos: 1.75801e+07 muA
** NormalTransistorNmos: 1.75791e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.18699e+06 muA


** Expected Voltages: 
** ibias: 1.16501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.95901  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.25  V
** outSourceVoltageBiasXXnXX1: 0.625  V
** outSourceVoltageBiasXXnXX2: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.09101  V
** innerStageBias: 0.590001  V
** innerTransistorStack1Load1: 4.08901  V
** out1: 3.21201  V
** sourceTransconductance: 1.94501  V
** inner: 0.625  V


.END