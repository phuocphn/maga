** Name: two_stage_single_output_op_amp_92_12

.MACRO two_stage_single_output_op_amp_92_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=42e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=550e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=168e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=256e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=15e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=65e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=65e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=65e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=42e-6
mMainBias12 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=20e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=550e-6
mTelescopicFirstStageLoad14 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=65e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=42e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=574e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=594e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mTelescopicFirstStageLoad19 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=256e-6
mMainBias20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=33e-6
mMainBias21 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=357e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.6001e-12
.EOM two_stage_single_output_op_amp_92_12

** Expected Performance Values: 
** Gain: 151 dB
** Power consumption: 4.28501 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 3.33701 MHz
** Transit frequency with error factor: 3.33504 MHz
** Slew rate: 9.96356 V/mu_s
** Phase margin: 61.8795°
** CMRR: 91 dB
** VoutMax: 4.61001 V
** VoutMin: 0.770001 V
** VcmMax: 4.51001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorNmos: 1.33431e+07 muA
** NormalTransistorNmos: 2.80221e+07 muA
** NormalTransistorPmos: -2.98219e+07 muA
** NormalTransistorPmos: -3.16809e+08 muA
** NormalTransistorNmos: 3.09511e+07 muA
** NormalTransistorNmos: 3.09511e+07 muA
** DiodeTransistorPmos: -3.09519e+07 muA
** NormalTransistorPmos: -3.09519e+07 muA
** NormalTransistorNmos: 3.78711e+08 muA
** NormalTransistorNmos: 3.09511e+07 muA
** NormalTransistorNmos: 3.09511e+07 muA
** NormalTransistorNmos: 3.97082e+08 muA
** DiodeTransistorNmos: 3.97081e+08 muA
** NormalTransistorPmos: -3.97081e+08 muA
** NormalTransistorPmos: -3.97082e+08 muA
** DiodeTransistorNmos: 2.98211e+07 muA
** NormalTransistorNmos: 2.98201e+07 muA
** DiodeTransistorNmos: 3.1681e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.33439e+07 muA
** DiodeTransistorPmos: -2.80229e+07 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.84401  V
** out: 2.5  V
** outFirstStage: 4.24201  V
** outInputVoltageBiasXXnXX1: 1.17801  V
** outSourceVoltageBiasXXnXX1: 0.589001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX1: 4.03901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.25201  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.79501  V
** inner: 0.589001  V


.END