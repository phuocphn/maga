** Name: two_stage_single_output_op_amp_175_2

.MACRO two_stage_single_output_op_amp_175_2 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=17e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=84e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=84e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=23e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
mSimpleFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=113e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=139e-6
mSecondStage1Transconductor9 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=557e-6
mSimpleFirstStageLoad10 outFirstStage outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=113e-6
mMainBias11 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=13e-6
mSimpleFirstStageStageBias12 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=205e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=84e-6
mSimpleFirstStageTransconductor14 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=349e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=139e-6
mSecondStage1StageBias16 out ibias sourcePmos sourcePmos pmos4 L=4e-6 W=600e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=84e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=349e-6
mMainBias19 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=25e-6
mMainBias20 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=159e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.1001e-12
.EOM two_stage_single_output_op_amp_175_2

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 6.81101 mW
** Area: 14981 (mu_m)^2
** Transit frequency: 3.47001 MHz
** Transit frequency with error factor: 3.44194 MHz
** Slew rate: 5.56318 V/mu_s
** Phase margin: 60.1606°
** CMRR: 88 dB
** VoutMax: 4.69001 V
** VoutMin: 0.300001 V
** VcmMax: 3.04001 V
** VcmMin: -0.0699999 V


** Expected Currents: 
** NormalTransistorNmos: 5.31791e+07 muA
** NormalTransistorPmos: -1.10519e+07 muA
** NormalTransistorPmos: -6.95419e+07 muA
** DiodeTransistorPmos: -4.26442e+08 muA
** NormalTransistorPmos: -4.26442e+08 muA
** NormalTransistorPmos: -4.26442e+08 muA
** DiodeTransistorPmos: -4.26442e+08 muA
** NormalTransistorNmos: 4.71564e+08 muA
** NormalTransistorNmos: 4.71564e+08 muA
** NormalTransistorPmos: -9.02429e+07 muA
** NormalTransistorPmos: -9.02439e+07 muA
** NormalTransistorPmos: -4.51209e+07 muA
** NormalTransistorPmos: -4.51209e+07 muA
** NormalTransistorNmos: 2.65258e+08 muA
** NormalTransistorNmos: 2.65257e+08 muA
** NormalTransistorPmos: -2.65257e+08 muA
** DiodeTransistorNmos: 1.10511e+07 muA
** DiodeTransistorNmos: 6.95411e+07 muA
** DiodeTransistorPmos: -5.31799e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.12301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX1: 0.727001  V
** outVoltageBiasXXnXX2: 0.899001  V
** outVoltageBiasXXpXX1: 3.84201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.68601  V
** innerStageBias: 4.67501  V
** innerTransistorStack1Load1: 3.68601  V
** out1: 2.37201  V
** sourceTransconductance: 3.31801  V
** innerTransconductance: 0.172001  V


.END