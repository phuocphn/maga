** Name: symmetrical_op_amp193

.MACRO symmetrical_op_amp193 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=10e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=86e-6
mSymmetricalFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=64e-6
mMainBias4 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=35e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=23e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=64e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=49e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias8 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=49e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=10e-6
mSymmetricalFirstStageTransconductor10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=75e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias11 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=5e-6 W=36e-6
mSecondStage1StageBias12 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=36e-6
mSymmetricalFirstStageTransconductor13 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=75e-6
mMainBias14 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=178e-6
mMainBias15 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=40e-6
mSymmetricalFirstStageLoad16 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=34e-6
mSymmetricalFirstStageLoad17 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=34e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=38e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor19 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=38e-6
mMainBias20 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=168e-6
mSymmetricalFirstStageLoad21 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=155e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor22 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=174e-6
mSecondStage1Transconductor23 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=174e-6
mSymmetricalFirstStageLoad24 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=155e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp193

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 3.23901 mW
** Area: 7734 (mu_m)^2
** Transit frequency: 3.54301 MHz
** Transit frequency with error factor: 3.54331 MHz
** Slew rate: 3.51957 V/mu_s
** Phase margin: 79.0682°
** CMRR: 142 dB
** negPSRR: 132 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 0.450001 V
** VcmMax: 4.81001 V
** VcmMin: 1.58001 V


** Expected Currents: 
** NormalTransistorNmos: 4.00041e+07 muA
** NormalTransistorNmos: 1.77684e+08 muA
** NormalTransistorPmos: -2.86751e+08 muA
** NormalTransistorPmos: -3.13919e+07 muA
** NormalTransistorPmos: -3.13929e+07 muA
** NormalTransistorPmos: -3.13919e+07 muA
** NormalTransistorPmos: -3.13929e+07 muA
** NormalTransistorNmos: 6.27821e+07 muA
** DiodeTransistorNmos: 6.27831e+07 muA
** NormalTransistorNmos: 3.13911e+07 muA
** NormalTransistorNmos: 3.13911e+07 muA
** NormalTransistorNmos: 3.52751e+07 muA
** NormalTransistorNmos: 3.52741e+07 muA
** NormalTransistorPmos: -3.52759e+07 muA
** NormalTransistorPmos: -3.52749e+07 muA
** NormalTransistorNmos: 3.52751e+07 muA
** NormalTransistorNmos: 3.52741e+07 muA
** NormalTransistorPmos: -3.52759e+07 muA
** NormalTransistorPmos: -3.52749e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 2.86752e+08 muA
** DiodeTransistorPmos: -4.00049e+07 muA
** DiodeTransistorPmos: -1.77683e+08 muA


** Expected Voltages: 
** ibias: 1.41901  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.851001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.611001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.711001  V
** outVoltageBiasXXpXX0: 3.99701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.93701  V
** innerStageBias: 0.206001  V
** innerTransconductance: 4.40001  V
** inner: 0.206001  V
** inner: 4.40001  V
** inner: 0.706001  V


.END