** Name: two_stage_single_output_op_amp_46_2

.MACRO two_stage_single_output_op_amp_46_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=64e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=201e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=7e-6 W=89e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=33e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=156e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=80e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=80e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=483e-6
mSecondStage1Transconductor10 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=389e-6
mFoldedCascodeFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=156e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=201e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=107e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=107e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=361e-6
mMainBias16 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=402e-6
mSecondStage1StageBias17 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad18 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=89e-6
mMainBias19 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=243e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.4001e-12
.EOM two_stage_single_output_op_amp_46_2

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 3.53501 mW
** Area: 14331 (mu_m)^2
** Transit frequency: 2.53701 MHz
** Transit frequency with error factor: 2.53664 MHz
** Slew rate: 5.20503 V/mu_s
** Phase margin: 60.1606°
** CMRR: 120 dB
** VoutMax: 4.82001 V
** VoutMin: 0.300001 V
** VcmMax: 3.80001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -7.50599e+07 muA
** NormalTransistorPmos: -1.21897e+08 muA
** NormalTransistorNmos: 9.66151e+07 muA
** NormalTransistorNmos: 1.52372e+08 muA
** NormalTransistorNmos: 9.66151e+07 muA
** NormalTransistorNmos: 1.52372e+08 muA
** DiodeTransistorPmos: -9.66159e+07 muA
** DiodeTransistorPmos: -9.66169e+07 muA
** NormalTransistorPmos: -9.66159e+07 muA
** NormalTransistorPmos: -9.66169e+07 muA
** NormalTransistorPmos: -1.11508e+08 muA
** NormalTransistorPmos: -5.57549e+07 muA
** NormalTransistorPmos: -5.57549e+07 muA
** NormalTransistorNmos: 1.85333e+08 muA
** NormalTransistorNmos: 1.85332e+08 muA
** NormalTransistorPmos: -1.85332e+08 muA
** DiodeTransistorNmos: 7.50591e+07 muA
** DiodeTransistorNmos: 1.21898e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX1: 0.926001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4  V
** innerTransistorStack2Load2: 3.99401  V
** out1: 2.78101  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.51401  V
** innerTransconductance: 0.371001  V


.END