** Name: two_stage_single_output_op_amp_55_11

.MACRO two_stage_single_output_op_amp_55_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=154e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=154e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias4 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=108e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=154e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=90e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=90e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=56e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mMainBias12 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=23e-6
mSecondStage1StageBias13 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=509e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=4e-6 W=154e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=62e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerOutputLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=201e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=363e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=363e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=593e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=555e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=201e-6
mMainBias22 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=241e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.7001e-12
.EOM two_stage_single_output_op_amp_55_11

** Expected Performance Values: 
** Gain: 175 dB
** Power consumption: 7.44401 mW
** Area: 14498 (mu_m)^2
** Transit frequency: 4.52201 MHz
** Transit frequency with error factor: 4.52235 MHz
** Slew rate: 3.92638 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 4.25 V
** VoutMin: 0.5 V
** VcmMax: 5.09001 V
** VcmMin: 0.800001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorNmos: 3.76311e+07 muA
** NormalTransistorPmos: -8.33149e+07 muA
** NormalTransistorPmos: -8.16329e+07 muA
** NormalTransistorPmos: -1.27444e+08 muA
** NormalTransistorPmos: -8.16329e+07 muA
** NormalTransistorPmos: -1.27444e+08 muA
** DiodeTransistorNmos: 8.16321e+07 muA
** NormalTransistorNmos: 8.16311e+07 muA
** NormalTransistorNmos: 8.16321e+07 muA
** DiodeTransistorNmos: 8.16311e+07 muA
** NormalTransistorNmos: 9.16231e+07 muA
** NormalTransistorNmos: 4.58111e+07 muA
** NormalTransistorNmos: 4.58111e+07 muA
** NormalTransistorNmos: 1.00151e+09 muA
** NormalTransistorNmos: 1.00151e+09 muA
** NormalTransistorPmos: -1.0015e+09 muA
** NormalTransistorPmos: -1.0015e+09 muA
** DiodeTransistorNmos: 8.33141e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -3.76319e+07 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.12401  V
** out: 2.5  V
** outFirstStage: 4.00301  V
** outVoltageBiasXXnXX1: 1.11001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.12601  V
** innerSourceLoad2: 0.563001  V
** innerTransistorStack1Load2: 0.562001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94001  V
** innerStageBias: 0.442001  V
** innerTransconductance: 4.56701  V


.END