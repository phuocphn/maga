** Name: two_stage_single_output_op_amp_58_10

.MACRO two_stage_single_output_op_amp_58_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=138e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=102e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=123e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=22e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=74e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=74e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=594e-6
mFoldedCascodeFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=22e-6
mMainBias12 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=82e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=142e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=142e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=123e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=587e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=333e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=102e-6
mMainBias21 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=529e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.5e-12
.EOM two_stage_single_output_op_amp_58_10

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 14.6931 mW
** Area: 5253 (mu_m)^2
** Transit frequency: 10.1301 MHz
** Transit frequency with error factor: 10.1181 MHz
** Slew rate: 9.47206 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** VoutMax: 4.25 V
** VoutMin: 0.170001 V
** VcmMax: 3.04001 V
** VcmMin: -0.389999 V


** Expected Currents: 
** NormalTransistorNmos: 2.03068e+08 muA
** NormalTransistorPmos: -5.31565e+08 muA
** NormalTransistorPmos: -3.38203e+08 muA
** NormalTransistorNmos: 1.18691e+08 muA
** NormalTransistorNmos: 1.81356e+08 muA
** NormalTransistorNmos: 1.18691e+08 muA
** NormalTransistorNmos: 1.81356e+08 muA
** DiodeTransistorPmos: -1.1869e+08 muA
** NormalTransistorPmos: -1.1869e+08 muA
** NormalTransistorPmos: -1.25326e+08 muA
** DiodeTransistorPmos: -1.25325e+08 muA
** NormalTransistorPmos: -6.26639e+07 muA
** NormalTransistorPmos: -6.26639e+07 muA
** NormalTransistorNmos: 1.48305e+09 muA
** NormalTransistorPmos: -1.48304e+09 muA
** NormalTransistorPmos: -1.48304e+09 muA
** DiodeTransistorNmos: 5.31566e+08 muA
** DiodeTransistorNmos: 3.38204e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -2.03067e+08 muA


** Expected Voltages: 
** ibias: 3.19701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.576001  V
** out: 2.5  V
** outFirstStage: 4.05901  V
** outSourceVoltageBiasXXpXX1: 4.10001  V
** outVoltageBiasXXnXX1: 1.13201  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.07401  V
** sourceGCC1: 0.371001  V
** sourceGCC2: 0.371001  V
** sourceTransconductance: 3.22101  V
** innerTransconductance: 4.62101  V
** inner: 4.09401  V


.END