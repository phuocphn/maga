** Name: two_stage_single_output_op_amp_115_9

.MACRO two_stage_single_output_op_amp_115_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=7e-6 W=27e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=537e-6
mMainBias4 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=22e-6
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=79e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=21e-6
mTelescopicFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=7e-6 W=144e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=30e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=30e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=30e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mMainBias13 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=7e-6 W=71e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=537e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=30e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=55e-6
mTelescopicFirstStageLoad17 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=79e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=529e-6
mTelescopicFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=9e-6 W=28e-6
mMainBias20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=27e-6
mMainBias21 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=26e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_115_9

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 5.58601 mW
** Area: 7656 (mu_m)^2
** Transit frequency: 3.83601 MHz
** Transit frequency with error factor: 3.83559 MHz
** Slew rate: 8.86421 V/mu_s
** Phase margin: 64.7443°
** CMRR: 135 dB
** VoutMax: 4.43001 V
** VoutMin: 0.700001 V
** VcmMax: 4.12001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 1.95291e+07 muA
** NormalTransistorPmos: -2.47619e+07 muA
** NormalTransistorPmos: -2.37079e+07 muA
** NormalTransistorNmos: 8.16401e+06 muA
** NormalTransistorNmos: 8.16301e+06 muA
** NormalTransistorPmos: -8.16499e+06 muA
** NormalTransistorPmos: -8.16399e+06 muA
** DiodeTransistorPmos: -8.16499e+06 muA
** NormalTransistorNmos: 4.00321e+07 muA
** NormalTransistorNmos: 4.00311e+07 muA
** NormalTransistorNmos: 8.16301e+06 muA
** NormalTransistorNmos: 8.16301e+06 muA
** NormalTransistorNmos: 1.02279e+09 muA
** DiodeTransistorNmos: 1.02279e+09 muA
** NormalTransistorPmos: -1.02278e+09 muA
** DiodeTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** DiodeTransistorNmos: 2.37071e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.95299e+07 muA


** Expected Voltages: 
** ibias: 1.13601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.88001  V
** out: 2.5  V
** outFirstStage: 3.86401  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX3: 0.556001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.24901  V
** innerStageBias: 0.485001  V
** out1: 3.30001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.555001  V


.END