** Name: two_stage_single_output_op_amp_74_5

.MACRO two_stage_single_output_op_amp_74_5 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=84e-6
mMainBias2 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=27e-6
mFoldedCascodeFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=70e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=7e-6 W=34e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=10e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=532e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=66e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=84e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=12e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=70e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=27e-6
mMainBias13 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=130e-6
mSecondStage1Transconductor14 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=171e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=4e-6 W=18e-6
mMainBias16 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=29e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=20e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=50e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=50e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=10e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=532e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=20e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_74_5

** Expected Performance Values: 
** Gain: 113 dB
** Power consumption: 3.56501 mW
** Area: 14669 (mu_m)^2
** Transit frequency: 3.04301 MHz
** Transit frequency with error factor: 3.04277 MHz
** Slew rate: 5.0673 V/mu_s
** Phase margin: 60.1606°
** CMRR: 126 dB
** VoutMax: 3.23001 V
** VoutMin: 0.590001 V
** VcmMax: 4.87001 V
** VcmMin: 1.52001 V


** Expected Currents: 
** NormalTransistorNmos: 1.07561e+07 muA
** NormalTransistorNmos: 4.79851e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorPmos: -3.56709e+07 muA
** NormalTransistorPmos: -2.28559e+07 muA
** NormalTransistorPmos: -3.56699e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28551e+07 muA
** DiodeTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.56261e+07 muA
** DiodeTransistorNmos: 2.56271e+07 muA
** NormalTransistorNmos: 1.28131e+07 muA
** NormalTransistorNmos: 1.28131e+07 muA
** NormalTransistorNmos: 5.72862e+08 muA
** NormalTransistorPmos: -5.72861e+08 muA
** DiodeTransistorPmos: -5.72862e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.07569e+07 muA
** NormalTransistorPmos: -1.07579e+07 muA
** DiodeTransistorPmos: -4.79859e+07 muA
** DiodeTransistorPmos: -4.79869e+07 muA


** Expected Voltages: 
** ibias: 1.22601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.59401  V
** out: 2.5  V
** outFirstStage: 0.999001  V
** outInputVoltageBiasXXpXX1: 2.66401  V
** outSourceVoltageBiasXXnXX1: 0.614001  V
** outSourceVoltageBiasXXpXX1: 3.83201  V
** outSourceVoltageBiasXXpXX2: 3.90501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** out1: 1.20401  V
** sourceGCC1: 3.82401  V
** sourceGCC2: 3.82401  V
** sourceTransconductance: 1.79701  V
** inner: 0.611001  V
** inner: 3.82601  V


.END