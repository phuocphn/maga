** Name: one_stage_single_output_op_amp73

.MACRO one_stage_single_output_op_amp73 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=56e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=6e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=12e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=228e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=71e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=56e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=61e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=61e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=74e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=100e-6
mFoldedCascodeFirstStageLoad12 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=3e-6 W=12e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=173e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=246e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=246e-6
mFoldedCascodeFirstStageLoad16 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=173e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp73

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 1.59901 mW
** Area: 2796 (mu_m)^2
** Transit frequency: 3.38701 MHz
** Transit frequency with error factor: 3.38683 MHz
** Slew rate: 3.50522 V/mu_s
** Phase margin: 88.8085°
** CMRR: 136 dB
** VoutMax: 4.13001 V
** VoutMin: 1.16001 V
** VcmMax: 5.25 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorNmos: 9.88751e+07 muA
** NormalTransistorPmos: -7.02609e+07 muA
** NormalTransistorPmos: -1.05497e+08 muA
** NormalTransistorPmos: -7.02609e+07 muA
** NormalTransistorPmos: -1.05497e+08 muA
** NormalTransistorNmos: 7.02601e+07 muA
** NormalTransistorNmos: 7.02601e+07 muA
** DiodeTransistorNmos: 7.02601e+07 muA
** NormalTransistorNmos: 7.04721e+07 muA
** NormalTransistorNmos: 7.04711e+07 muA
** NormalTransistorNmos: 3.52361e+07 muA
** NormalTransistorNmos: 3.52361e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.88759e+07 muA
** DiodeTransistorPmos: -9.8875e+07 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.28101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.702001  V
** innerStageBias: 0.606001  V
** out1: 1.56101  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.92901  V


.END