** Name: two_stage_single_output_op_amp_161_1

.MACRO two_stage_single_output_op_amp_161_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=18e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=52e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=29e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=567e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=567e-6
mSimpleFirstStageLoad8 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=244e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=386e-6
mSimpleFirstStageLoad10 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=244e-6
mMainBias11 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=64e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=71e-6
mSimpleFirstStageStageBias13 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSimpleFirstStageTransconductor14 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=11e-6
mSimpleFirstStageLoad15 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=52e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=7e-6 W=124e-6
mSecondStage1StageBias17 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=342e-6
mSimpleFirstStageLoad18 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=29e-6
mSimpleFirstStageTransconductor19 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=11e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_161_1

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 5.54901 mW
** Area: 11978 (mu_m)^2
** Transit frequency: 2.74901 MHz
** Transit frequency with error factor: 2.74712 MHz
** Slew rate: 3.50014 V/mu_s
** Phase margin: 77.3494°
** CMRR: 118 dB
** VoutMax: 4.71001 V
** VoutMin: 0.350001 V
** VcmMax: 3.16001 V
** VcmMin: -0.179999 V


** Expected Currents: 
** NormalTransistorNmos: 3.05291e+07 muA
** NormalTransistorNmos: 3.39571e+07 muA
** NormalTransistorPmos: -2.61908e+08 muA
** NormalTransistorPmos: -2.61908e+08 muA
** DiodeTransistorPmos: -2.61908e+08 muA
** NormalTransistorNmos: 2.69981e+08 muA
** NormalTransistorNmos: 2.69982e+08 muA
** NormalTransistorNmos: 2.69981e+08 muA
** NormalTransistorNmos: 2.69982e+08 muA
** NormalTransistorPmos: -1.61449e+07 muA
** NormalTransistorPmos: -1.61459e+07 muA
** NormalTransistorPmos: -8.07199e+06 muA
** NormalTransistorPmos: -8.07199e+06 muA
** NormalTransistorNmos: 4.95382e+08 muA
** NormalTransistorPmos: -4.95381e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -3.05299e+07 muA
** DiodeTransistorPmos: -3.39579e+07 muA


** Expected Voltages: 
** ibias: 1.12201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.755001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 3.79101  V
** outVoltageBiasXXpXX2: 4.15001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.58001  V
** innerTransistorStack1Load2: 0.488001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.488001  V
** out1: 2.40801  V
** sourceTransconductance: 3.26601  V


.END