** Name: two_stage_single_output_op_amp_114_7

.MACRO two_stage_single_output_op_amp_114_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=7e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=117e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=8e-6
mTelescopicFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=10e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=10e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias11 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=19e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
mTelescopicFirstStageStageBias14 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=117e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=549e-6
mTelescopicFirstStageLoad16 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mMainBias17 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=6e-6
mMainBias18 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=67e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.5e-12
.EOM two_stage_single_output_op_amp_114_7

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 2.12701 mW
** Area: 5846 (mu_m)^2
** Transit frequency: 7.33301 MHz
** Transit frequency with error factor: 7.32758 MHz
** Slew rate: 11.1137 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** VoutMax: 4.83001 V
** VoutMin: 0.170001 V
** VcmMax: 4.51001 V
** VcmMin: 1.52001 V


** Expected Currents: 
** NormalTransistorNmos: 9.06101e+06 muA
** NormalTransistorPmos: -6.80099e+06 muA
** NormalTransistorPmos: -7.54319e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorNmos: 1.13525e+08 muA
** DiodeTransistorNmos: 1.13524e+08 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 2.86032e+08 muA
** NormalTransistorPmos: -2.86031e+08 muA
** DiodeTransistorNmos: 6.80001e+06 muA
** NormalTransistorNmos: 6.79901e+06 muA
** DiodeTransistorNmos: 7.54311e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.06199e+06 muA


** Expected Voltages: 
** ibias: 0.572001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4  V
** out: 2.5  V
** outFirstStage: 4.26501  V
** outInputVoltageBiasXXnXX1: 1.37401  V
** outSourceVoltageBiasXXnXX1: 0.687001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.25901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.685001  V


.END