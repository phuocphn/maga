** Name: two_stage_single_output_op_amp_81_11

.MACRO two_stage_single_output_op_amp_81_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=17e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=17e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=5e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=88e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=302e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=16e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=545e-6
mSecondStage1StageBias13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=563e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=6e-6 W=17e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=300e-6
mMainBias16 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=45e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=126e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=212e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=212e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=432e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=420e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=126e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.10001e-12
.EOM two_stage_single_output_op_amp_81_11

** Expected Performance Values: 
** Gain: 177 dB
** Power consumption: 4.75001 mW
** Area: 9810 (mu_m)^2
** Transit frequency: 4.22001 MHz
** Transit frequency with error factor: 4.21955 MHz
** Slew rate: 4.00455 V/mu_s
** Phase margin: 60.1606°
** CMRR: 142 dB
** VoutMax: 4.28001 V
** VoutMin: 0.710001 V
** VcmMax: 5.20001 V
** VcmMin: 1.33001 V


** Expected Currents: 
** NormalTransistorNmos: 2.97833e+08 muA
** NormalTransistorNmos: 4.41441e+07 muA
** NormalTransistorPmos: -2.06009e+07 muA
** NormalTransistorPmos: -3.08999e+07 muA
** NormalTransistorPmos: -2.06049e+07 muA
** NormalTransistorPmos: -3.09059e+07 muA
** DiodeTransistorNmos: 2.06021e+07 muA
** NormalTransistorNmos: 2.06031e+07 muA
** NormalTransistorNmos: 2.06041e+07 muA
** DiodeTransistorNmos: 2.06031e+07 muA
** NormalTransistorNmos: 2.06001e+07 muA
** NormalTransistorNmos: 2.06011e+07 muA
** NormalTransistorNmos: 1.03001e+07 muA
** NormalTransistorNmos: 1.03001e+07 muA
** NormalTransistorNmos: 5.36153e+08 muA
** NormalTransistorNmos: 5.36152e+08 muA
** NormalTransistorPmos: -5.36152e+08 muA
** NormalTransistorPmos: -5.36153e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.97832e+08 muA
** DiodeTransistorPmos: -4.41449e+07 muA


** Expected Voltages: 
** ibias: 1.18001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.17201  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.23401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.672001  V
** innerStageBias: 0.554001  V
** innerTransistorStack1Load2: 0.670001  V
** out1: 1.36901  V
** sourceGCC1: 4.41501  V
** sourceGCC2: 4.41501  V
** sourceTransconductance: 1.94401  V
** innerStageBias: 0.625  V
** innerTransconductance: 4.71101  V


.END