** Name: two_stage_single_output_op_amp_29_7

.MACRO two_stage_single_output_op_amp_29_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=118e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=275e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mSimpleFirstStageStageBias5 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=273e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=14e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=129e-6
mSecondStage1StageBias8 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=299e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=14e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=48e-6
mMainBias11 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=262e-6
mSecondStage1Transconductor12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=275e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_29_7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 7.88101 mW
** Area: 3072 (mu_m)^2
** Transit frequency: 6.19601 MHz
** Transit frequency with error factor: 6.15674 MHz
** Slew rate: 10.1922 V/mu_s
** Phase margin: 60.1606°
** CMRR: 88 dB
** negPSRR: 130 dB
** posPSRR: 86 dB
** VoutMax: 4.83001 V
** VoutMin: 0.150001 V
** VcmMax: 4.68001 V
** VcmMin: 1.87001 V


** Expected Currents: 
** NormalTransistorNmos: 4.79401e+07 muA
** NormalTransistorPmos: -9.5041e+08 muA
** DiodeTransistorPmos: -1.3467e+08 muA
** NormalTransistorPmos: -1.3467e+08 muA
** NormalTransistorNmos: 2.6934e+08 muA
** NormalTransistorNmos: 2.69339e+08 muA
** NormalTransistorNmos: 1.34671e+08 muA
** NormalTransistorNmos: 1.34671e+08 muA
** NormalTransistorNmos: 2.98439e+08 muA
** NormalTransistorPmos: -2.98438e+08 muA
** DiodeTransistorNmos: 9.50411e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.79409e+07 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.715001  V
** out: 2.5  V
** outFirstStage: 4.27001  V
** outVoltageBiasXXpXX0: 3.98401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.153001  V
** out1: 4.27001  V
** sourceTransconductance: 1.34501  V


.END