** Name: two_stage_single_output_op_amp_45_9

.MACRO two_stage_single_output_op_amp_45_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=49e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=71e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=358e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=71e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=51e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
mMainBias7 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=44e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=22e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=22e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=49e-6
mMainBias12 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=26e-6
mSecondStage1StageBias13 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=358e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=51e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=79e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=79e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=102e-6
mMainBias19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=480e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=496e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=192e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=9e-6 W=284e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_45_9

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 6.89501 mW
** Area: 9426 (mu_m)^2
** Transit frequency: 5.65001 MHz
** Transit frequency with error factor: 5.64971 MHz
** Slew rate: 6.08342 V/mu_s
** Phase margin: 62.4525°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.760001 V
** VcmMax: 4.02001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.96371e+07 muA
** NormalTransistorPmos: -1.30119e+08 muA
** NormalTransistorPmos: -1.35229e+08 muA
** NormalTransistorNmos: 2.78601e+07 muA
** NormalTransistorNmos: 4.19021e+07 muA
** NormalTransistorNmos: 2.78601e+07 muA
** NormalTransistorNmos: 4.19021e+07 muA
** DiodeTransistorPmos: -2.78609e+07 muA
** NormalTransistorPmos: -2.78609e+07 muA
** NormalTransistorPmos: -2.78609e+07 muA
** NormalTransistorPmos: -2.80809e+07 muA
** NormalTransistorPmos: -1.40409e+07 muA
** NormalTransistorPmos: -1.40409e+07 muA
** NormalTransistorNmos: 9.60252e+08 muA
** DiodeTransistorNmos: 9.60251e+08 muA
** NormalTransistorPmos: -9.60251e+08 muA
** DiodeTransistorNmos: 1.3012e+08 muA
** NormalTransistorNmos: 1.30121e+08 muA
** DiodeTransistorNmos: 1.3523e+08 muA
** DiodeTransistorNmos: 1.3523e+08 muA
** DiodeTransistorPmos: -4.96379e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.16601  V
** inputVoltageBiasXXnXX2: 1.11001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.583001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.47201  V
** out1: 4.26101  V
** sourceGCC1: 0.551001  V
** sourceGCC2: 0.551001  V
** sourceTransconductance: 3.23601  V
** inner: 0.584001  V


.END