** Name: two_stage_single_output_op_amp_205_12

.MACRO two_stage_single_output_op_amp_205_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=40e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=40e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=8e-6
mMainBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=18e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=254e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias7 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=121e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=178e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=40e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=187e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=58e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=18e-6
mMainBias14 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=276e-6
mSecondStage1StageBias15 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=254e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=40e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=187e-6
mMainBias18 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=216e-6
mSimpleFirstStageLoad19 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=216e-6
mSimpleFirstStageLoad20 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=216e-6
mSimpleFirstStageLoad21 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=521e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=557e-6
mMainBias23 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=69e-6
mSecondStage1Transconductor24 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad25 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=521e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.4001e-12
.EOM two_stage_single_output_op_amp_205_12

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 12.7691 mW
** Area: 12720 (mu_m)^2
** Transit frequency: 7.15201 MHz
** Transit frequency with error factor: 7.14923 MHz
** Slew rate: 6.74075 V/mu_s
** Phase margin: 60.1606°
** CMRR: 111 dB
** VoutMax: 4.25 V
** VoutMin: 1.68001 V
** VcmMax: 4.72001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 1.42147e+08 muA
** NormalTransistorNmos: 1.80501e+08 muA
** NormalTransistorPmos: -1.04086e+08 muA
** DiodeTransistorNmos: 2.65816e+08 muA
** NormalTransistorNmos: 2.65817e+08 muA
** NormalTransistorNmos: 2.65816e+08 muA
** DiodeTransistorNmos: 2.65817e+08 muA
** NormalTransistorPmos: -3.25176e+08 muA
** NormalTransistorPmos: -3.25177e+08 muA
** NormalTransistorPmos: -3.25176e+08 muA
** NormalTransistorPmos: -3.25177e+08 muA
** NormalTransistorNmos: 1.18722e+08 muA
** NormalTransistorNmos: 1.18721e+08 muA
** NormalTransistorNmos: 5.93611e+07 muA
** NormalTransistorNmos: 5.93611e+07 muA
** NormalTransistorNmos: 1.46669e+09 muA
** DiodeTransistorNmos: 1.46669e+09 muA
** NormalTransistorPmos: -1.46668e+09 muA
** NormalTransistorPmos: -1.46668e+09 muA
** DiodeTransistorNmos: 1.04087e+08 muA
** NormalTransistorNmos: 1.04086e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.42146e+08 muA
** DiodeTransistorPmos: -1.805e+08 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.08401  V
** inputVoltageBiasXXpXX2: 3.93401  V
** out: 2.5  V
** outFirstStage: 4.05401  V
** outSourceVoltageBiasXXnXX1: 1.04201  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15001  V
** innerStageBias: 0.498001  V
** innerTransistorStack1Load1: 1.15001  V
** innerTransistorStack1Load2: 4.43601  V
** innerTransistorStack2Load2: 4.43601  V
** out1: 2.11801  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.61801  V
** inner: 1.03601  V


.END