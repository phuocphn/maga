** Name: two_stage_single_output_op_amp_87_1

.MACRO two_stage_single_output_op_amp_87_1 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=83e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=105e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=27e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=9e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=6e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=83e-6
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=519e-6
mTelescopicFirstStageLoad8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=73e-6
mMainBias9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mTelescopicFirstStageLoad10 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=6e-6 W=11e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=49e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=49e-6
mMainBias13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=100e-6
mSecondStage1StageBias14 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=445e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=6e-6 W=11e-6
mMainBias16 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=24e-6
mTelescopicFirstStageStageBias17 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=51e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.90001e-12
.EOM two_stage_single_output_op_amp_87_1

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 3.61201 mW
** Area: 5855 (mu_m)^2
** Transit frequency: 7.08401 MHz
** Transit frequency with error factor: 7.08432 MHz
** Slew rate: 9.74487 V/mu_s
** Phase margin: 60.1606°
** CMRR: 141 dB
** VoutMax: 4.57001 V
** VoutMin: 0.150001 V
** VcmMax: 3.85001 V
** VcmMin: 0.920001 V


** Expected Currents: 
** NormalTransistorNmos: 1.79981e+07 muA
** NormalTransistorPmos: -2.70219e+07 muA
** NormalTransistorPmos: -1.13329e+08 muA
** NormalTransistorPmos: -1.99009e+07 muA
** NormalTransistorPmos: -1.99009e+07 muA
** DiodeTransistorNmos: 1.99001e+07 muA
** NormalTransistorNmos: 1.99001e+07 muA
** NormalTransistorNmos: 1.99001e+07 muA
** NormalTransistorPmos: -5.77979e+07 muA
** NormalTransistorPmos: -1.98999e+07 muA
** NormalTransistorPmos: -1.98999e+07 muA
** NormalTransistorNmos: 5.04321e+08 muA
** NormalTransistorPmos: -5.0432e+08 muA
** DiodeTransistorNmos: 2.70211e+07 muA
** DiodeTransistorNmos: 1.1333e+08 muA
** DiodeTransistorPmos: -1.79989e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.00201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.556001  V
** outVoltageBiasXXnXX0: 0.558001  V
** outVoltageBiasXXpXX1: 1.64301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21401  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 2.99001  V
** sourceGCC2: 2.99001  V


.END