** Name: two_stage_single_output_op_amp_151_9

.MACRO two_stage_single_output_op_amp_151_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=11e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=11e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=5e-6
mMainBias4 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=221e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=44e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=11e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=95e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=221e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=11e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=44e-6
mSimpleFirstStageLoad14 FirstStageYinnerOutputLoad1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=301e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=134e-6
mMainBias16 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=266e-6
mSimpleFirstStageLoad18 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=301e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.80001e-12
.EOM two_stage_single_output_op_amp_151_9

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 14.9981 mW
** Area: 2628 (mu_m)^2
** Transit frequency: 11.2771 MHz
** Transit frequency with error factor: 11.2501 MHz
** Slew rate: 10.6281 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 1.46001 V
** VcmMax: 5.25 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorPmos: -5.88629e+07 muA
** NormalTransistorPmos: -7.02799e+06 muA
** DiodeTransistorNmos: 8.79581e+07 muA
** NormalTransistorNmos: 8.79591e+07 muA
** NormalTransistorNmos: 8.79601e+07 muA
** DiodeTransistorNmos: 8.79591e+07 muA
** NormalTransistorPmos: -1.2986e+08 muA
** NormalTransistorPmos: -1.2986e+08 muA
** NormalTransistorNmos: 8.38031e+07 muA
** NormalTransistorNmos: 4.19021e+07 muA
** NormalTransistorNmos: 4.19021e+07 muA
** NormalTransistorNmos: 2.65403e+09 muA
** DiodeTransistorNmos: 2.65403e+09 muA
** NormalTransistorPmos: -2.65402e+09 muA
** DiodeTransistorNmos: 5.88621e+07 muA
** NormalTransistorNmos: 5.88611e+07 muA
** DiodeTransistorNmos: 7.02701e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.87001  V
** inputVoltageBiasXXnXX2: 0.581001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.935001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack1Load1: 1.15601  V
** sourceTransconductance: 1.94501  V
** inner: 0.935001  V


.END