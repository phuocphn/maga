** Name: two_stage_single_output_op_amp_47_12

.MACRO two_stage_single_output_op_amp_47_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=8e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=241e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=54e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=72e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=72e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=241e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=54e-6
mMainBias13 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=449e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=283e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=283e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=339e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=339e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=468e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=478e-6
mMainBias21 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=48e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=449e-6
mMainBias24 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=44e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.2001e-12
.EOM two_stage_single_output_op_amp_47_12

** Expected Performance Values: 
** Gain: 151 dB
** Power consumption: 14.9681 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 8.43301 MHz
** Transit frequency with error factor: 8.43228 MHz
** Slew rate: 33.2405 V/mu_s
** Phase margin: 60.1606°
** CMRR: 122 dB
** VoutMax: 4.25 V
** VoutMin: 1.85001 V
** VcmMax: 3.48001 V
** VcmMin: -0.0799999 V


** Expected Currents: 
** NormalTransistorNmos: 9.97361e+07 muA
** NormalTransistorPmos: -4.48209e+07 muA
** NormalTransistorPmos: -4.88829e+07 muA
** NormalTransistorNmos: 4.76854e+08 muA
** NormalTransistorNmos: 7.15279e+08 muA
** NormalTransistorNmos: 4.76856e+08 muA
** NormalTransistorNmos: 7.15281e+08 muA
** NormalTransistorPmos: -4.76853e+08 muA
** NormalTransistorPmos: -4.76854e+08 muA
** NormalTransistorPmos: -4.76855e+08 muA
** NormalTransistorPmos: -4.76854e+08 muA
** NormalTransistorPmos: -4.76851e+08 muA
** NormalTransistorPmos: -2.38425e+08 muA
** NormalTransistorPmos: -2.38425e+08 muA
** NormalTransistorNmos: 1.34956e+09 muA
** DiodeTransistorNmos: 1.34956e+09 muA
** NormalTransistorPmos: -1.34955e+09 muA
** NormalTransistorPmos: -1.34955e+09 muA
** DiodeTransistorNmos: 4.48201e+07 muA
** NormalTransistorNmos: 4.48191e+07 muA
** DiodeTransistorNmos: 4.88821e+07 muA
** DiodeTransistorNmos: 4.88811e+07 muA
** DiodeTransistorPmos: -9.97369e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.10001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.77201  V
** out: 2.5  V
** outFirstStage: 4.03901  V
** outInputVoltageBiasXXnXX1: 2.25801  V
** outSourceVoltageBiasXXnXX1: 1.12901  V
** outSourceVoltageBiasXXnXX2: 0.888001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.12901  V
** innerTransistorStack1Load2: 4.49301  V
** innerTransistorStack2Load2: 4.49301  V
** sourceGCC1: 0.908001  V
** sourceGCC2: 0.908001  V
** sourceTransconductance: 3.68901  V
** innerTransconductance: 4.60301  V
** inner: 1.12201  V


.END