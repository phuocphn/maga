** Name: two_stage_single_output_op_amp_203_7

.MACRO two_stage_single_output_op_amp_203_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=6e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
mMainBias4 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=58e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=105e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=28e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=38e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=19e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=281e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=6e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=38e-6
mSimpleFirstStageLoad13 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=590e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=570e-6
mMainBias15 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=385e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=253e-6
mSimpleFirstStageLoad17 outFirstStage ibias sourcePmos sourcePmos pmos4 L=5e-6 W=590e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_203_7

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 2.02701 mW
** Area: 13336 (mu_m)^2
** Transit frequency: 3.94201 MHz
** Transit frequency with error factor: 3.92085 MHz
** Slew rate: 3.71497 V/mu_s
** Phase margin: 60.1606°
** CMRR: 95 dB
** VoutMax: 4.80001 V
** VoutMin: 0.150001 V
** VcmMax: 5.24001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorPmos: -5.53449e+07 muA
** NormalTransistorPmos: -3.69469e+07 muA
** DiodeTransistorNmos: 4.79771e+07 muA
** NormalTransistorNmos: 4.79781e+07 muA
** NormalTransistorNmos: 4.79791e+07 muA
** DiodeTransistorNmos: 4.79781e+07 muA
** NormalTransistorPmos: -5.70249e+07 muA
** NormalTransistorPmos: -5.70249e+07 muA
** NormalTransistorNmos: 1.80941e+07 muA
** NormalTransistorNmos: 1.80931e+07 muA
** NormalTransistorNmos: 9.04701e+06 muA
** NormalTransistorNmos: 9.04701e+06 muA
** NormalTransistorNmos: 1.78998e+08 muA
** NormalTransistorPmos: -1.78997e+08 muA
** DiodeTransistorNmos: 5.53441e+07 muA
** DiodeTransistorNmos: 3.69461e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.710001  V
** inputVoltageBiasXXnXX2: 0.556001  V
** out: 2.5  V
** outFirstStage: 4.23701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.155001  V
** innerTransistorStack1Load1: 1.15601  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V


.END