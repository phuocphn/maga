** Name: two_stage_single_output_op_amp_30_7

.MACRO two_stage_single_output_op_amp_30_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=35e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=266e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=288e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=228e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=16e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=266e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=35e-6
mMainBias9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=57e-6
mSecondStage1StageBias10 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=328e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=16e-6
mSecondStage1Transconductor12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=288e-6
mMainBias14 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=158e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_30_7

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 3.08701 mW
** Area: 5137 (mu_m)^2
** Transit frequency: 5.89801 MHz
** Transit frequency with error factor: 5.86088 MHz
** Slew rate: 9.23146 V/mu_s
** Phase margin: 60.1606°
** CMRR: 88 dB
** negPSRR: 133 dB
** posPSRR: 87 dB
** VoutMax: 4.84001 V
** VoutMin: 0.170001 V
** VcmMax: 4.68001 V
** VcmMin: 1.93001 V


** Expected Currents: 
** NormalTransistorNmos: 4.75041e+07 muA
** NormalTransistorPmos: -3.31059e+07 muA
** DiodeTransistorPmos: -1.28257e+08 muA
** NormalTransistorPmos: -1.28257e+08 muA
** NormalTransistorNmos: 2.56514e+08 muA
** DiodeTransistorNmos: 2.56513e+08 muA
** NormalTransistorNmos: 1.28258e+08 muA
** NormalTransistorNmos: 1.28258e+08 muA
** NormalTransistorNmos: 2.70367e+08 muA
** NormalTransistorPmos: -2.70366e+08 muA
** DiodeTransistorNmos: 3.31051e+07 muA
** NormalTransistorNmos: 3.31051e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.75049e+07 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.28301  V
** out: 2.5  V
** outFirstStage: 4.27801  V
** outInputVoltageBiasXXnXX1: 1.17801  V
** outSourceVoltageBiasXXnXX1: 0.589001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.27801  V
** sourceTransconductance: 1.34501  V
** inner: 0.589001  V


.END