** Name: two_stage_single_output_op_amp_12_9

.MACRO two_stage_single_output_op_amp_12_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=19e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=66e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=24e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=15e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=19e-6
mMainBias9 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=16e-6
mSecondStage1StageBias10 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=66e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=15e-6
mMainBias12 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mSimpleFirstStageLoad13 FirstStageYinnerSourceLoad1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=9e-6 W=217e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=14e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=14e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=317e-6
mSimpleFirstStageLoad17 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=9e-6 W=217e-6
mMainBias18 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=32e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_12_9

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 3.78601 mW
** Area: 6834 (mu_m)^2
** Transit frequency: 2.94901 MHz
** Transit frequency with error factor: 2.9466 MHz
** Slew rate: 4.31995 V/mu_s
** Phase margin: 64.1713°
** CMRR: 94 dB
** negPSRR: 94 dB
** posPSRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 1.01001 V
** VcmMax: 4.81001 V
** VcmMin: 0.840001 V


** Expected Currents: 
** NormalTransistorNmos: 2.81161e+07 muA
** NormalTransistorNmos: 2.68171e+07 muA
** NormalTransistorPmos: -1.48137e+08 muA
** NormalTransistorPmos: -9.85799e+06 muA
** NormalTransistorPmos: -9.85899e+06 muA
** NormalTransistorPmos: -9.85799e+06 muA
** NormalTransistorPmos: -9.85899e+06 muA
** NormalTransistorNmos: 1.97151e+07 muA
** NormalTransistorNmos: 9.85701e+06 muA
** NormalTransistorNmos: 9.85701e+06 muA
** NormalTransistorNmos: 5.24337e+08 muA
** DiodeTransistorNmos: 5.24336e+08 muA
** NormalTransistorPmos: -5.24336e+08 muA
** DiodeTransistorNmos: 1.48138e+08 muA
** NormalTransistorNmos: 1.48137e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.81169e+07 muA
** DiodeTransistorPmos: -2.68179e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.68801  V
** outInputVoltageBiasXXnXX1: 1.42001  V
** outSourceVoltageBiasXXnXX1: 0.710001  V
** outVoltageBiasXXpXX0: 3.71301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.83801  V
** innerTransistorStack1Load1: 4.40101  V
** innerTransistorStack2Load1: 4.40101  V
** sourceTransconductance: 1.86101  V
** inner: 0.710001  V


.END