** Name: two_stage_single_output_op_amp_55_9

.MACRO two_stage_single_output_op_amp_55_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=29e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=29e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=6e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=270e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=20e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=23e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=22e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=10e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=75e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=270e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=4e-6 W=29e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerOutputLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=128e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=64e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=64e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=246e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=128e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=39e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=14e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_55_9

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 4.60301 mW
** Area: 6995 (mu_m)^2
** Transit frequency: 3.56101 MHz
** Transit frequency with error factor: 3.56051 MHz
** Slew rate: 3.81196 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 4.25 V
** VoutMin: 1.33001 V
** VcmMax: 5.13001 V
** VcmMin: 0.810001 V


** Expected Currents: 
** NormalTransistorPmos: -1.80039e+07 muA
** NormalTransistorPmos: -6.46299e+06 muA
** NormalTransistorPmos: -1.73279e+07 muA
** NormalTransistorPmos: -2.95459e+07 muA
** NormalTransistorPmos: -1.73279e+07 muA
** NormalTransistorPmos: -2.95459e+07 muA
** DiodeTransistorNmos: 1.73271e+07 muA
** NormalTransistorNmos: 1.73261e+07 muA
** NormalTransistorNmos: 1.73271e+07 muA
** DiodeTransistorNmos: 1.73261e+07 muA
** NormalTransistorNmos: 2.44331e+07 muA
** NormalTransistorNmos: 1.22171e+07 muA
** NormalTransistorNmos: 1.22171e+07 muA
** NormalTransistorNmos: 8.17123e+08 muA
** DiodeTransistorNmos: 8.17122e+08 muA
** NormalTransistorPmos: -8.17122e+08 muA
** DiodeTransistorNmos: 1.80031e+07 muA
** NormalTransistorNmos: 1.80021e+07 muA
** DiodeTransistorNmos: 6.46201e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.73201  V
** outSourceVoltageBiasXXnXX1: 0.866001  V
** outSourceVoltageBiasXXpXX1: 4.15901  V
** outVoltageBiasXXnXX2: 0.569001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.22901  V
** innerSourceLoad2: 0.656001  V
** innerTransistorStack1Load2: 0.656001  V
** sourceGCC1: 4.03801  V
** sourceGCC2: 4.03801  V
** sourceTransconductance: 1.85401  V
** inner: 0.864001  V


.END