** Name: symmetrical_op_amp9

.MACRO symmetrical_op_amp9 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=39e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSymmetricalFirstStageLoad4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=39e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=63e-6
mMainBias6 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=8e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=90e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=90e-6
mMainBias9 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=33e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=4e-6 W=70e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=70e-6
mSymmetricalFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=5e-6 W=189e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=125e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias14 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=125e-6
mMainBias15 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=5e-6 W=61e-6
mSymmetricalFirstStageTransconductor16 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=81e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias17 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=4e-6 W=32e-6
mMainBias18 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=15e-6
mSecondStage1StageBias19 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=4e-6 W=40e-6
mSymmetricalFirstStageTransconductor20 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=81e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp9

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 0.762001 mW
** Area: 5626 (mu_m)^2
** Transit frequency: 2.72001 MHz
** Transit frequency with error factor: 2.71971 MHz
** Slew rate: 3.50045 V/mu_s
** Phase margin: 74.4846°
** CMRR: 146 dB
** negPSRR: 52 dB
** posPSRR: 88 dB
** VoutMax: 4.31001 V
** VoutMin: 0.300001 V
** VcmMax: 4.02001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 1.99091e+07 muA
** NormalTransistorPmos: -2.40999e+06 muA
** NormalTransistorPmos: -9.75899e+06 muA
** DiodeTransistorNmos: 1.51881e+07 muA
** DiodeTransistorNmos: 1.51881e+07 muA
** NormalTransistorPmos: -3.03769e+07 muA
** NormalTransistorPmos: -1.51889e+07 muA
** NormalTransistorPmos: -1.51889e+07 muA
** NormalTransistorNmos: 3.50451e+07 muA
** NormalTransistorNmos: 3.50441e+07 muA
** NormalTransistorPmos: -3.50459e+07 muA
** NormalTransistorPmos: -3.50469e+07 muA
** NormalTransistorPmos: -3.48329e+07 muA
** NormalTransistorPmos: -3.48339e+07 muA
** NormalTransistorNmos: 3.48321e+07 muA
** NormalTransistorNmos: 3.48311e+07 muA
** DiodeTransistorNmos: 2.40901e+06 muA
** DiodeTransistorNmos: 9.75801e+06 muA
** DiodeTransistorPmos: -1.99099e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.22501  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 3.68601  V
** inOutputTransconductanceComplementarySecondStage: 0.710001  V
** inSourceTransconductanceComplementarySecondStage: 0.556001  V
** innerComplementarySecondStage: 4.18501  V
** inputVoltageBiasXXnXX0: 0.573001  V
** out: 2.5  V
** outFirstStage: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.26801  V
** innerStageBias: 4.69101  V
** innerTransconductance: 0.151001  V
** inner: 4.74201  V
** inner: 0.151001  V


.END