** Name: two_stage_single_output_op_amp_3_5

.MACRO two_stage_single_output_op_amp_3_5 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=131e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=17e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=39e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=9e-6 W=11e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=131e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=131e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=471e-6
mSimpleFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=64e-6
mMainBias10 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=46e-6
mSimpleFirstStageTransconductor11 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=15e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=98e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=11e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=38e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=9e-6 W=131e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=15e-6
mMainBias17 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.5e-12
.EOM two_stage_single_output_op_amp_3_5

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 1.53301 mW
** Area: 8818 (mu_m)^2
** Transit frequency: 3.84601 MHz
** Transit frequency with error factor: 3.83078 MHz
** Slew rate: 5.00166 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** negPSRR: 94 dB
** posPSRR: 203 dB
** VoutMax: 3.03001 V
** VoutMin: 0.150001 V
** VcmMax: 3.36001 V
** VcmMin: 0.210001 V


** Expected Currents: 
** NormalTransistorNmos: 1.07471e+07 muA
** NormalTransistorPmos: -9.16999e+06 muA
** NormalTransistorPmos: -3.85189e+07 muA
** DiodeTransistorNmos: 4.99281e+07 muA
** NormalTransistorNmos: 4.99271e+07 muA
** NormalTransistorNmos: 4.99281e+07 muA
** NormalTransistorPmos: -9.98529e+07 muA
** NormalTransistorPmos: -4.99269e+07 muA
** NormalTransistorPmos: -4.99269e+07 muA
** NormalTransistorNmos: 1.28215e+08 muA
** NormalTransistorPmos: -1.28214e+08 muA
** DiodeTransistorPmos: -1.28215e+08 muA
** DiodeTransistorNmos: 9.16901e+06 muA
** DiodeTransistorNmos: 3.85181e+07 muA
** DiodeTransistorPmos: -1.07479e+07 muA
** NormalTransistorPmos: -1.07489e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.10001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.769001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.46201  V
** outSourceVoltageBiasXXpXX1: 3.73101  V
** outVoltageBiasXXnXX0: 0.571001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.80801  V
** inner: 3.72401  V


.END