** Name: two_stage_single_output_op_amp_88_3

.MACRO two_stage_single_output_op_amp_88_3 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=27e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=9e-6 W=27e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=51e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=250e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=27e-6
mMainBias8 inputVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=373e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=292e-6
mTelescopicFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=27e-6
mMainBias11 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=378e-6
mTelescopicFirstStageLoad12 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=47e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=75e-6
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=75e-6
mSecondStage1StageBias15 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=438e-6
mMainBias16 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=20e-6
mSecondStage1StageBias17 out inputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=599e-6
mTelescopicFirstStageLoad18 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=47e-6
mTelescopicFirstStageStageBias19 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=160e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_88_3

** Expected Performance Values: 
** Gain: 150 dB
** Power consumption: 3.97001 mW
** Area: 14991 (mu_m)^2
** Transit frequency: 2.51501 MHz
** Transit frequency with error factor: 2.51527 MHz
** Slew rate: 17.7984 V/mu_s
** Phase margin: 68.182°
** CMRR: 131 dB
** VoutMax: 4.31001 V
** VoutMin: 0.300001 V
** VcmMax: 3.94001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorNmos: 1.51593e+08 muA
** NormalTransistorNmos: 1.50381e+08 muA
** NormalTransistorPmos: -2.01559e+07 muA
** NormalTransistorPmos: -5.71499e+06 muA
** NormalTransistorPmos: -5.71499e+06 muA
** DiodeTransistorNmos: 5.71401e+06 muA
** DiodeTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorPmos: -1.63025e+08 muA
** NormalTransistorPmos: -5.71599e+06 muA
** NormalTransistorPmos: -5.71599e+06 muA
** NormalTransistorNmos: 4.40517e+08 muA
** NormalTransistorPmos: -4.40516e+08 muA
** NormalTransistorPmos: -4.40517e+08 muA
** DiodeTransistorNmos: 2.01551e+07 muA
** DiodeTransistorPmos: -1.51592e+08 muA
** DiodeTransistorPmos: -1.5038e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.10001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.611001  V
** inputVoltageBiasXXpXX2: 1.93601  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outVoltageBiasXXpXX1: 2.29101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.22401  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 3.02001  V
** sourceGCC2: 3.02001  V
** innerStageBias: 2.85001  V


.END