** Name: symmetrical_op_amp24

.MACRO symmetrical_op_amp24 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias4 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSymmetricalFirstStageLoad5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=522e-6
mSymmetricalFirstStageLoad6 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=522e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias9 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos4 L=3e-6 W=14e-6
mSymmetricalFirstStageTransconductor10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=37e-6
mSecondStage1StageBias11 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=85e-6
mSymmetricalFirstStageTransconductor12 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=37e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=493e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=493e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=248e-6
mSecondStage1Transconductor16 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=248e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp24

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 5.45901 mW
** Area: 5096 (mu_m)^2
** Transit frequency: 13.8731 MHz
** Transit frequency with error factor: 13.8726 MHz
** Slew rate: 26.2294 V/mu_s
** Phase margin: 74.4846°
** CMRR: 144 dB
** negPSRR: 49 dB
** posPSRR: 41 dB
** VoutMax: 4.49001 V
** VoutMin: 1.15001 V
** VcmMax: 4.67001 V
** VcmMin: 0.880001 V


** Expected Currents: 
** NormalTransistorNmos: 1.25361e+07 muA
** DiodeTransistorPmos: -2.73967e+08 muA
** DiodeTransistorPmos: -2.73967e+08 muA
** NormalTransistorNmos: 5.47934e+08 muA
** NormalTransistorNmos: 2.73968e+08 muA
** NormalTransistorNmos: 2.73968e+08 muA
** NormalTransistorNmos: 2.63265e+08 muA
** NormalTransistorNmos: 2.63264e+08 muA
** NormalTransistorPmos: -2.63264e+08 muA
** NormalTransistorPmos: -2.63263e+08 muA
** DiodeTransistorNmos: 2.58162e+08 muA
** DiodeTransistorNmos: 2.58163e+08 muA
** NormalTransistorPmos: -2.58161e+08 muA
** NormalTransistorPmos: -2.58162e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.25369e+07 muA


** Expected Voltages: 
** ibias: 0.584001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.90401  V
** inSourceStageBiasComplementarySecondStage: 0.960001  V
** inSourceTransconductanceComplementarySecondStage: 4.26401  V
** innerComplementarySecondStage: 1.91501  V
** out: 2.5  V
** outFirstStage: 4.26401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.79801  V
** innerStageBias: 1.31801  V
** innerTransconductance: 4.81101  V
** inner: 4.80801  V


.END