** Name: two_stage_single_output_op_amp_47_7

.MACRO two_stage_single_output_op_amp_47_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=52e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=90e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=56e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=141e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=141e-6
mMainBias8 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=21e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=589e-6
mFoldedCascodeFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=56e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=196e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=111e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=111e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=273e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=273e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=586e-6
mMainBias17 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=360e-6
mMainBias18 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=297e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=196e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12e-12
.EOM two_stage_single_output_op_amp_47_7

** Expected Performance Values: 
** Gain: 134 dB
** Power consumption: 3.31701 mW
** Area: 14981 (mu_m)^2
** Transit frequency: 5.30401 MHz
** Transit frequency with error factor: 5.30445 MHz
** Slew rate: 4.66774 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.81001 V
** VoutMin: 0.150001 V
** VcmMax: 4.08001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.34671e+07 muA
** NormalTransistorPmos: -4.04329e+07 muA
** NormalTransistorPmos: -3.30149e+07 muA
** NormalTransistorNmos: 5.63421e+07 muA
** NormalTransistorNmos: 8.95181e+07 muA
** NormalTransistorNmos: 5.63421e+07 muA
** NormalTransistorNmos: 8.95181e+07 muA
** NormalTransistorPmos: -5.63429e+07 muA
** NormalTransistorPmos: -5.63439e+07 muA
** NormalTransistorPmos: -5.63429e+07 muA
** NormalTransistorPmos: -5.63439e+07 muA
** NormalTransistorPmos: -6.63489e+07 muA
** NormalTransistorPmos: -3.31749e+07 muA
** NormalTransistorPmos: -3.31749e+07 muA
** NormalTransistorNmos: 3.77366e+08 muA
** NormalTransistorPmos: -3.77365e+08 muA
** DiodeTransistorNmos: 4.04321e+07 muA
** DiodeTransistorNmos: 3.30141e+07 muA
** DiodeTransistorPmos: -1.34679e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.943001  V
** inputVoltageBiasXXnXX2: 0.555001  V
** inputVoltageBiasXXpXX1: 3.88501  V
** out: 2.5  V
** outFirstStage: 4.24801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.26701  V
** innerTransistorStack1Load2: 4.62801  V
** innerTransistorStack2Load2: 4.62801  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.22901  V


.END