** Name: symmetrical_op_amp146

.MACRO symmetrical_op_amp146 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias3 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=496e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=82e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=82e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=163e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=163e-6
mSymmetricalFirstStageLoad9 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=53e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=4e-6 W=92e-6
mSecondStage1Transconductor11 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=92e-6
mSymmetricalFirstStageLoad12 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=53e-6
mSymmetricalFirstStageStageBias13 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=309e-6
mSymmetricalFirstStageStageBias14 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=155e-6
mSymmetricalFirstStageTransconductor15 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=592e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias16 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=496e-6
mSecondStage1StageBias17 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=1e-6 W=163e-6
mSymmetricalFirstStageTransconductor18 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=592e-6
mMainBias19 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp146

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 4.89801 mW
** Area: 11426 (mu_m)^2
** Transit frequency: 16.5791 MHz
** Transit frequency with error factor: 16.5795 MHz
** Slew rate: 30.958 V/mu_s
** Phase margin: 74.4846°
** CMRR: 142 dB
** negPSRR: 40 dB
** posPSRR: 63 dB
** VoutMax: 3.84001 V
** VoutMin: 0.550001 V
** VcmMax: 3 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.53459e+07 muA
** NormalTransistorNmos: 1.56645e+08 muA
** NormalTransistorNmos: 1.56644e+08 muA
** NormalTransistorNmos: 1.56645e+08 muA
** NormalTransistorNmos: 1.56644e+08 muA
** NormalTransistorPmos: -3.13288e+08 muA
** NormalTransistorPmos: -3.13287e+08 muA
** NormalTransistorPmos: -1.56644e+08 muA
** NormalTransistorPmos: -1.56644e+08 muA
** NormalTransistorNmos: 3.10456e+08 muA
** NormalTransistorNmos: 3.10455e+08 muA
** NormalTransistorPmos: -3.10455e+08 muA
** DiodeTransistorPmos: -3.10456e+08 muA
** NormalTransistorPmos: -3.10455e+08 muA
** NormalTransistorNmos: 3.10456e+08 muA
** NormalTransistorNmos: 3.10455e+08 muA
** DiodeTransistorNmos: 2.53451e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** inStageBiasComplementarySecondStage: 4.17101  V
** innerComplementarySecondStage: 3.27901  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.953001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.29701  V
** innerTransistorStack1Load1: 0.173001  V
** innerTransistorStack2Load1: 0.173001  V
** sourceTransconductance: 3.36101  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END