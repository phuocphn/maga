** Name: two_stage_single_output_op_amp_65_1

.MACRO two_stage_single_output_op_amp_65_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=7e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=5e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=88e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=88e-6
mMainBias8 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=117e-6
mFoldedCascodeFirstStageLoad10 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=21e-6
mMainBias11 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=41e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=33e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=33e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=190e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=68e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=68e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=5e-6 W=478e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=495e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=190e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_65_1

** Expected Performance Values: 
** Gain: 113 dB
** Power consumption: 3.03101 mW
** Area: 8428 (mu_m)^2
** Transit frequency: 3.40401 MHz
** Transit frequency with error factor: 3.4039 MHz
** Slew rate: 8.40224 V/mu_s
** Phase margin: 62.4525°
** CMRR: 131 dB
** VoutMax: 4.68001 V
** VoutMin: 0.580001 V
** VcmMax: 3 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.00071e+07 muA
** NormalTransistorNmos: 4.67001e+06 muA
** NormalTransistorNmos: 3.81501e+07 muA
** NormalTransistorNmos: 5.75511e+07 muA
** NormalTransistorNmos: 3.81501e+07 muA
** NormalTransistorNmos: 5.75511e+07 muA
** NormalTransistorPmos: -3.81509e+07 muA
** NormalTransistorPmos: -3.81519e+07 muA
** NormalTransistorPmos: -3.81509e+07 muA
** NormalTransistorPmos: -3.81519e+07 muA
** NormalTransistorPmos: -3.88049e+07 muA
** NormalTransistorPmos: -3.88059e+07 muA
** NormalTransistorPmos: -1.94019e+07 muA
** NormalTransistorPmos: -1.94019e+07 muA
** NormalTransistorNmos: 4.66387e+08 muA
** NormalTransistorPmos: -4.66386e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.00079e+07 muA
** DiodeTransistorPmos: -4.67099e+06 muA


** Expected Voltages: 
** ibias: 1.18701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.982001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX2: 4.11201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40001  V
** innerTransistorStack1Load2: 4.48601  V
** innerTransistorStack2Load2: 4.48601  V
** out1: 4.18101  V
** sourceGCC1: 0.527001  V
** sourceGCC2: 0.527001  V
** sourceTransconductance: 3.46201  V


.END