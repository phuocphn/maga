** Name: two_stage_single_output_op_amp_71_6

.MACRO two_stage_single_output_op_amp_71_6 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=93e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mSecondStage1StageBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=11e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=12e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=593e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=193e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=337e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=337e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=112e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=591e-6
mMainBias13 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=100e-6
mSecondStage1Transconductor14 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=588e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=93e-6
mMainBias16 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerLoad2 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=439e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=593e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=439e-6
mMainBias23 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.8001e-12
.EOM two_stage_single_output_op_amp_71_6

** Expected Performance Values: 
** Gain: 148 dB
** Power consumption: 11.7331 mW
** Area: 8406 (mu_m)^2
** Transit frequency: 14.2611 MHz
** Transit frequency with error factor: 14.2516 MHz
** Slew rate: 11.1391 V/mu_s
** Phase margin: 60.1606°
** CMRR: 110 dB
** VoutMax: 3.78001 V
** VoutMin: 0.300001 V
** VcmMax: 4.66001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 2.30961e+07 muA
** NormalTransistorNmos: 1.11687e+08 muA
** NormalTransistorPmos: -5.07669e+08 muA
** NormalTransistorPmos: -1.77318e+08 muA
** NormalTransistorPmos: -2.84294e+08 muA
** NormalTransistorPmos: -1.77318e+08 muA
** NormalTransistorPmos: -2.84294e+08 muA
** DiodeTransistorNmos: 1.77319e+08 muA
** NormalTransistorNmos: 1.77319e+08 muA
** NormalTransistorNmos: 2.13954e+08 muA
** NormalTransistorNmos: 2.13953e+08 muA
** NormalTransistorNmos: 1.06978e+08 muA
** NormalTransistorNmos: 1.06978e+08 muA
** NormalTransistorNmos: 1.12564e+09 muA
** NormalTransistorNmos: 1.12564e+09 muA
** NormalTransistorPmos: -1.12563e+09 muA
** DiodeTransistorPmos: -1.12563e+09 muA
** DiodeTransistorNmos: 5.0767e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.30969e+07 muA
** NormalTransistorPmos: -2.30979e+07 muA
** DiodeTransistorPmos: -1.11686e+08 muA
** DiodeTransistorPmos: -1.11686e+08 muA


** Expected Voltages: 
** ibias: 0.567001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.21801  V
** outSourceVoltageBiasXXpXX1: 4.10901  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX1: 0.917001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.555001  V
** innerStageBias: 0.362001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 0.361001  V
** inner: 4.10901  V


.END