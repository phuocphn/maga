** Name: two_stage_single_output_op_amp_77_5

.MACRO two_stage_single_output_op_amp_77_5 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=7e-6 W=30e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=68e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=4e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=3e-6 W=35e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=28e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=266e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=35e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=50e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=68e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=50e-6
mMainBias14 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=247e-6
mSecondStage1Transconductor15 out outFirstStage sourceNmos sourceNmos nmos4 L=10e-6 W=285e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=30e-6
mMainBias17 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=178e-6
mFoldedCascodeFirstStageLoad18 FirstStageYinnerOutputLoad2 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=138e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=9e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=9e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=28e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=266e-6
mFoldedCascodeFirstStageLoad23 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=138e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_77_5

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 5.33301 mW
** Area: 9306 (mu_m)^2
** Transit frequency: 4.07401 MHz
** Transit frequency with error factor: 4.07396 MHz
** Slew rate: 3.99929 V/mu_s
** Phase margin: 60.7336°
** CMRR: 142 dB
** VoutMax: 3.02001 V
** VoutMin: 0.580001 V
** VcmMax: 4.66001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 8.47561e+07 muA
** NormalTransistorNmos: 1.18456e+08 muA
** NormalTransistorPmos: -1.85569e+07 muA
** NormalTransistorPmos: -3.04599e+07 muA
** NormalTransistorPmos: -1.85569e+07 muA
** NormalTransistorPmos: -3.04599e+07 muA
** DiodeTransistorNmos: 1.85561e+07 muA
** DiodeTransistorNmos: 1.85551e+07 muA
** NormalTransistorNmos: 1.85561e+07 muA
** NormalTransistorNmos: 1.85551e+07 muA
** NormalTransistorNmos: 2.38081e+07 muA
** NormalTransistorNmos: 2.38081e+07 muA
** NormalTransistorNmos: 1.19041e+07 muA
** NormalTransistorNmos: 1.19041e+07 muA
** NormalTransistorNmos: 7.92494e+08 muA
** NormalTransistorPmos: -7.92493e+08 muA
** DiodeTransistorPmos: -7.92494e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -8.47569e+07 muA
** NormalTransistorPmos: -8.47579e+07 muA
** DiodeTransistorPmos: -1.18455e+08 muA
** DiodeTransistorPmos: -1.18455e+08 muA


** Expected Voltages: 
** ibias: 1.30201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.981001  V
** outInputVoltageBiasXXpXX1: 2.45201  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.72601  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.18601  V
** innerStageBias: 0.747001  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.554001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.89401  V
** inner: 3.72601  V


.END