** Name: two_stage_single_output_op_amp_15_2

.MACRO two_stage_single_output_op_amp_15_2 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSecondStage1StageBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=33e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSecondStage1Transconductor6 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=261e-6
mMainBias7 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mSecondStage1Transconductor8 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=72e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=52e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=12e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=3e-6 W=25e-6
mMainBias13 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=9e-6
mSecondStage1StageBias14 out ibias sourcePmos sourcePmos pmos4 L=7e-6 W=383e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=12e-6
mMainBias16 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=104e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_15_2

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 1.00201 mW
** Area: 6469 (mu_m)^2
** Transit frequency: 2.90401 MHz
** Transit frequency with error factor: 2.89884 MHz
** Slew rate: 3.50003 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** negPSRR: 98 dB
** posPSRR: 131 dB
** VoutMax: 4.65001 V
** VoutMin: 0.390001 V
** VcmMax: 3.01001 V
** VcmMin: 0.0300001 V


** Expected Currents: 
** NormalTransistorNmos: 1.15331e+07 muA
** NormalTransistorPmos: -2.77799e+06 muA
** NormalTransistorPmos: -3.21049e+07 muA
** DiodeTransistorNmos: 7.88701e+06 muA
** NormalTransistorNmos: 7.88701e+06 muA
** NormalTransistorPmos: -1.57769e+07 muA
** NormalTransistorPmos: -1.57779e+07 muA
** NormalTransistorPmos: -7.88799e+06 muA
** NormalTransistorPmos: -7.88799e+06 muA
** NormalTransistorNmos: 1.18233e+08 muA
** NormalTransistorNmos: 1.18232e+08 muA
** NormalTransistorPmos: -1.18232e+08 muA
** DiodeTransistorNmos: 2.77701e+06 muA
** DiodeTransistorNmos: 3.21041e+07 muA
** DiodeTransistorPmos: -1.15339e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.09001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.586001  V
** inputVoltageBiasXXpXX1: 3.73701  V
** out: 2.5  V
** outFirstStage: 0.598001  V
** outVoltageBiasXXnXX1: 0.794001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.625  V
** out1: 0.598001  V
** sourceTransconductance: 3.25501  V
** innerTransconductance: 0.193001  V


.END