** Name: two_stage_single_output_op_amp_22_5

.MACRO two_stage_single_output_op_amp_22_5 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=66e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=8e-6 W=66e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=34e-6
mMainBias4 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=2e-6 W=26e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=567e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=173e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=517e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=66e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=66e-6
mMainBias11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=138e-6
mSimpleFirstStageTransconductor12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=37e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=173e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=567e-6
mMainBias15 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=26e-6
mSecondStage1StageBias16 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=517e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=37e-6
mMainBias18 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=65e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_22_5

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 1.91601 mW
** Area: 9966 (mu_m)^2
** Transit frequency: 2.70301 MHz
** Transit frequency with error factor: 2.69742 MHz
** Slew rate: 6.92813 V/mu_s
** Phase margin: 61.3065°
** CMRR: 98 dB
** negPSRR: 92 dB
** posPSRR: 95 dB
** VoutMax: 4.02001 V
** VoutMin: 0.350001 V
** VcmMax: 3.12001 V
** VcmMin: 0.550001 V


** Expected Currents: 
** NormalTransistorNmos: 1.04477e+08 muA
** NormalTransistorPmos: -2.53799e+07 muA
** DiodeTransistorNmos: 1.57141e+07 muA
** DiodeTransistorNmos: 1.57141e+07 muA
** NormalTransistorNmos: 1.57141e+07 muA
** NormalTransistorNmos: 1.57141e+07 muA
** NormalTransistorPmos: -3.14309e+07 muA
** DiodeTransistorPmos: -3.14319e+07 muA
** NormalTransistorPmos: -1.57149e+07 muA
** NormalTransistorPmos: -1.57149e+07 muA
** NormalTransistorNmos: 2.01873e+08 muA
** NormalTransistorPmos: -2.01872e+08 muA
** DiodeTransistorPmos: -2.01871e+08 muA
** DiodeTransistorNmos: 2.53791e+07 muA
** DiodeTransistorPmos: -1.04476e+08 muA
** NormalTransistorPmos: -1.04477e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.45401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.756001  V
** outInputVoltageBiasXXpXX1: 3.52201  V
** outSourceVoltageBiasXXpXX1: 4.26101  V
** outSourceVoltageBiasXXpXX2: 4.22801  V
** outVoltageBiasXXnXX0: 0.568001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.555001  V
** out1: 1.11001  V
** sourceTransconductance: 3.47001  V
** inner: 4.26101  V
** inner: 4.22501  V


.END