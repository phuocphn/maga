** Name: two_stage_single_output_op_amp_124_10

.MACRO two_stage_single_output_op_amp_124_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=39e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=98e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=5e-6
mTelescopicFirstStageLoad5 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=295e-6
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=295e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=10e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad9 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=29e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=131e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=9e-6 W=131e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=39e-6
mMainBias13 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mSecondStage1StageBias14 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=460e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=29e-6
mMainBias16 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mTelescopicFirstStageStageBias17 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=98e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=295e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=238e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=567e-6
mTelescopicFirstStageLoad21 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=5e-6 W=295e-6
mMainBias22 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=17e-6
mMainBias23 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=11e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.2001e-12
.EOM two_stage_single_output_op_amp_124_10

** Expected Performance Values: 
** Gain: 150 dB
** Power consumption: 5.94201 mW
** Area: 14985 (mu_m)^2
** Transit frequency: 3.04701 MHz
** Transit frequency with error factor: 3.04725 MHz
** Slew rate: 3.84872 V/mu_s
** Phase margin: 60.1606°
** CMRR: 153 dB
** VoutMax: 4.46001 V
** VoutMin: 0.220001 V
** VcmMax: 3.80001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 1.71111e+07 muA
** NormalTransistorNmos: 6.03953e+08 muA
** NormalTransistorPmos: -2.91909e+07 muA
** NormalTransistorPmos: -1.88589e+07 muA
** NormalTransistorNmos: 2.77221e+07 muA
** NormalTransistorNmos: 2.77221e+07 muA
** DiodeTransistorPmos: -2.77229e+07 muA
** NormalTransistorPmos: -2.77239e+07 muA
** NormalTransistorPmos: -2.77229e+07 muA
** DiodeTransistorPmos: -2.77239e+07 muA
** NormalTransistorNmos: 7.43031e+07 muA
** DiodeTransistorNmos: 7.43021e+07 muA
** NormalTransistorNmos: 2.77231e+07 muA
** NormalTransistorNmos: 2.77231e+07 muA
** NormalTransistorNmos: 4.53863e+08 muA
** NormalTransistorPmos: -4.53862e+08 muA
** NormalTransistorPmos: -4.53863e+08 muA
** DiodeTransistorNmos: 2.91901e+07 muA
** NormalTransistorNmos: 2.91901e+07 muA
** DiodeTransistorNmos: 1.88581e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.71119e+07 muA
** DiodeTransistorPmos: -6.03952e+08 muA


** Expected Voltages: 
** ibias: 0.622001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.50401  V
** out: 2.5  V
** outFirstStage: 4.10801  V
** outInputVoltageBiasXXnXX1: 1.18801  V
** outSourceVoltageBiasXXnXX1: 0.594001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX1: 2.58901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerOutputLoad2: 3.54801  V
** innerSourceLoad2: 4.27401  V
** innerTransistorStack1Load2: 4.27401  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 3.36401  V
** inner: 0.594001  V


.END