** Name: two_stage_single_output_op_amp_9_12

.MACRO two_stage_single_output_op_amp_9_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=18e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=87e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=310e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=123e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=38e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=86e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=6e-6 W=197e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=87e-6
mMainBias10 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=67e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=310e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=86e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=555e-6
mSimpleFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=123e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=405e-6
mSecondStage1Transconductor16 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=221e-6
mMainBias18 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=359e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.6001e-12
.EOM two_stage_single_output_op_amp_9_12

** Expected Performance Values: 
** Gain: 142 dB
** Power consumption: 10.2071 mW
** Area: 9492 (mu_m)^2
** Transit frequency: 7.38301 MHz
** Transit frequency with error factor: 7.37917 MHz
** Slew rate: 6.95817 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** negPSRR: 112 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 0.840001 V
** VcmMax: 4.45001 V
** VcmMin: 0.75 V


** Expected Currents: 
** NormalTransistorNmos: 3.69481e+07 muA
** NormalTransistorNmos: 3.04602e+08 muA
** NormalTransistorPmos: -3.43356e+08 muA
** NormalTransistorPmos: -5.46009e+07 muA
** NormalTransistorPmos: -5.46009e+07 muA
** DiodeTransistorPmos: -5.46009e+07 muA
** NormalTransistorNmos: 1.092e+08 muA
** NormalTransistorNmos: 5.46001e+07 muA
** NormalTransistorNmos: 5.46001e+07 muA
** NormalTransistorNmos: 1.2373e+09 muA
** DiodeTransistorNmos: 1.2373e+09 muA
** NormalTransistorPmos: -1.23729e+09 muA
** NormalTransistorPmos: -1.23729e+09 muA
** DiodeTransistorNmos: 3.43357e+08 muA
** NormalTransistorNmos: 3.43357e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.69489e+07 muA
** DiodeTransistorPmos: -3.04601e+08 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.03401  V
** out: 2.5  V
** outFirstStage: 4.02401  V
** outInputVoltageBiasXXnXX1: 1.24401  V
** outSourceVoltageBiasXXnXX1: 0.622001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.21401  V
** out1: 3.48401  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.58801  V
** inner: 0.622001  V


.END