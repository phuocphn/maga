** Name: two_stage_single_output_op_amp_160_4

.MACRO two_stage_single_output_op_amp_160_4 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=45e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=13e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=235e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=13e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=108e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=73e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=203e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=107e-6
mSecondStage1Transconductor10 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=432e-6
mSimpleFirstStageLoad11 outFirstStage outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=203e-6
mMainBias12 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=340e-6
mSimpleFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=235e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=73e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=203e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=108e-6
mSecondStage1StageBias18 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=132e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=4e-6 W=312e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=340e-6
mMainBias21 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=85e-6
mMainBias22 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16e-12
.EOM two_stage_single_output_op_amp_160_4

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 10.5051 mW
** Area: 14902 (mu_m)^2
** Transit frequency: 2.69601 MHz
** Transit frequency with error factor: 2.65105 MHz
** Slew rate: 3.82489 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 3.91001 V
** VoutMin: 0.300001 V
** VcmMax: 3.03001 V
** VcmMin: -0.0799999 V


** Expected Currents: 
** NormalTransistorNmos: 9.14371e+07 muA
** NormalTransistorPmos: -8.61789e+07 muA
** NormalTransistorPmos: -5.16829e+07 muA
** NormalTransistorPmos: -7.91965e+08 muA
** NormalTransistorPmos: -7.91964e+08 muA
** DiodeTransistorPmos: -7.91965e+08 muA
** NormalTransistorNmos: 8.22935e+08 muA
** NormalTransistorNmos: 8.22935e+08 muA
** NormalTransistorPmos: -6.19389e+07 muA
** DiodeTransistorPmos: -6.19399e+07 muA
** NormalTransistorPmos: -3.09689e+07 muA
** NormalTransistorPmos: -3.09689e+07 muA
** NormalTransistorNmos: 2.05818e+08 muA
** NormalTransistorNmos: 2.05817e+08 muA
** NormalTransistorPmos: -2.05817e+08 muA
** NormalTransistorPmos: -2.05816e+08 muA
** DiodeTransistorNmos: 8.61781e+07 muA
** DiodeTransistorNmos: 5.16821e+07 muA
** DiodeTransistorPmos: -9.14379e+07 muA
** NormalTransistorPmos: -9.14389e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.42701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.25401  V
** outSourceVoltageBiasXXpXX1: 4.12701  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX1: 0.705001  V
** outVoltageBiasXXnXX2: 0.892001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.68601  V
** out1: 2.37201  V
** sourceTransconductance: 3.28901  V
** innerStageBias: 4.28501  V
** innerTransconductance: 0.150001  V
** inner: 4.125  V


.END