** Name: one_stage_single_output_op_amp55

.MACRO one_stage_single_output_op_amp55 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=37e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=37e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=20e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=165e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=37e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=72e-6
mFoldedCascodeFirstStageLoad10 out FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=3e-6 W=37e-6
mMainBias11 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=69e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerOutputLoad2 outInputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=276e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=222e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=222e-6
mFoldedCascodeFirstStageLoad15 out outInputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=276e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp55

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 2.57001 mW
** Area: 2105 (mu_m)^2
** Transit frequency: 5.96001 MHz
** Transit frequency with error factor: 5.96037 MHz
** Slew rate: 5.58349 V/mu_s
** Phase margin: 87.6626°
** CMRR: 138 dB
** VoutMax: 4.07001 V
** VoutMin: 1.06001 V
** VcmMax: 5.19001 V
** VcmMin: 0.810001 V


** Expected Currents: 
** NormalTransistorNmos: 1.37674e+08 muA
** NormalTransistorPmos: -1.12092e+08 muA
** NormalTransistorPmos: -1.83132e+08 muA
** NormalTransistorPmos: -1.12092e+08 muA
** NormalTransistorPmos: -1.83132e+08 muA
** DiodeTransistorNmos: 1.12093e+08 muA
** NormalTransistorNmos: 1.12092e+08 muA
** NormalTransistorNmos: 1.12093e+08 muA
** DiodeTransistorNmos: 1.12092e+08 muA
** NormalTransistorNmos: 1.4208e+08 muA
** NormalTransistorNmos: 7.10391e+07 muA
** NormalTransistorNmos: 7.10391e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.37673e+08 muA
** DiodeTransistorPmos: -1.37672e+08 muA


** Expected Voltages: 
** ibias: 0.622001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outInputVoltageBiasXXpXX1: 3.03601  V
** outSourceVoltageBiasXXpXX1: 4.22101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.46401  V
** innerSourceLoad2: 0.732001  V
** innerTransistorStack1Load2: 0.730001  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.90601  V


.END