** Name: two_stage_single_output_op_amp_44_3

.MACRO two_stage_single_output_op_amp_44_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=12e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=146e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=8e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=41e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=100e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=100e-6
mMainBias9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=41e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=67e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=41e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=54e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=146e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=50e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=435e-6
mSecondStage1StageBias18 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=596e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=8e-6 W=128e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.80001e-12
.EOM two_stage_single_output_op_amp_44_3

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 2.94501 mW
** Area: 7491 (mu_m)^2
** Transit frequency: 2.66101 MHz
** Transit frequency with error factor: 2.66074 MHz
** Slew rate: 5.55608 V/mu_s
** Phase margin: 60.1606°
** CMRR: 129 dB
** VoutMax: 4.45001 V
** VoutMin: 0.520001 V
** VcmMax: 3.88001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.70741e+07 muA
** NormalTransistorNmos: 3.55831e+07 muA
** NormalTransistorNmos: 4.35551e+07 muA
** NormalTransistorNmos: 6.53991e+07 muA
** NormalTransistorNmos: 4.35551e+07 muA
** NormalTransistorNmos: 6.53991e+07 muA
** NormalTransistorPmos: -4.35559e+07 muA
** NormalTransistorPmos: -4.35559e+07 muA
** DiodeTransistorPmos: -4.35559e+07 muA
** NormalTransistorPmos: -4.36909e+07 muA
** NormalTransistorPmos: -2.18449e+07 muA
** NormalTransistorPmos: -2.18449e+07 muA
** NormalTransistorNmos: 3.85465e+08 muA
** NormalTransistorPmos: -3.85464e+08 muA
** NormalTransistorPmos: -3.85465e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.70749e+07 muA
** DiodeTransistorPmos: -3.55839e+07 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.929001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX2: 4.21401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.04701  V
** out1: 3.09101  V
** sourceGCC1: 0.534001  V
** sourceGCC2: 0.534001  V
** sourceTransconductance: 3.39601  V
** innerStageBias: 4.57801  V


.END