** Name: two_stage_single_output_op_amp_196_11

.MACRO two_stage_single_output_op_amp_196_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=85e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=124e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=9e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=40e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=40e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=11e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=15e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=85e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=54e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=40e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=509e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=40e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=528e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=124e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=54e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=37e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mSimpleFirstStageLoad19 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=599e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=592e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=528e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=599e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=17e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.80001e-12
.EOM two_stage_single_output_op_amp_196_11

** Expected Performance Values: 
** Gain: 106 dB
** Power consumption: 14.9791 mW
** Area: 14539 (mu_m)^2
** Transit frequency: 4.54901 MHz
** Transit frequency with error factor: 4.38382 MHz
** Slew rate: 4.28764 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.29001 V
** VoutMin: 0.710001 V
** VcmMax: 4.66001 V
** VcmMin: 1.56001 V


** Expected Currents: 
** NormalTransistorNmos: 3.70291e+07 muA
** NormalTransistorNmos: 3.00231e+07 muA
** NormalTransistorPmos: -3.44289e+07 muA
** DiodeTransistorNmos: 1.17359e+09 muA
** DiodeTransistorNmos: 1.17359e+09 muA
** NormalTransistorNmos: 1.17359e+09 muA
** NormalTransistorNmos: 1.17359e+09 muA
** NormalTransistorPmos: -1.19072e+09 muA
** NormalTransistorPmos: -1.19072e+09 muA
** NormalTransistorNmos: 3.42831e+07 muA
** DiodeTransistorNmos: 3.42821e+07 muA
** NormalTransistorNmos: 1.71421e+07 muA
** NormalTransistorNmos: 1.71421e+07 muA
** NormalTransistorNmos: 5.02823e+08 muA
** NormalTransistorNmos: 5.02822e+08 muA
** NormalTransistorPmos: -5.02822e+08 muA
** NormalTransistorPmos: -5.02823e+08 muA
** DiodeTransistorNmos: 3.44281e+07 muA
** NormalTransistorNmos: 3.44271e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.70299e+07 muA
** DiodeTransistorPmos: -3.00239e+07 muA


** Expected Voltages: 
** ibias: 1.125  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.12701  V
** outInputVoltageBiasXXnXX1: 1.41201  V
** outSourceVoltageBiasXXnXX1: 0.706001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 3.68701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.10801  V
** innerTransistorStack2Load1: 1.10801  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.570001  V
** innerTransconductance: 4.64801  V
** inner: 0.703001  V


.END