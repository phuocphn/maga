** Name: two_stage_single_output_op_amp_40_10

.MACRO two_stage_single_output_op_amp_40_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=177e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=202e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=241e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=5e-6 W=241e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=578e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=66e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=56e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=202e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=177e-6
mMainBias11 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=100e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=599e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=56e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=338e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=241e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=371e-6
mSecondStage1Transconductor17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad18 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=241e-6
mMainBias19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=267e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.3001e-12
.EOM two_stage_single_output_op_amp_40_10

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 11.2741 mW
** Area: 14931 (mu_m)^2
** Transit frequency: 6.50701 MHz
** Transit frequency with error factor: 6.50416 MHz
** Slew rate: 6.13304 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** negPSRR: 115 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 0.260001 V
** VcmMax: 3.87001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 1.97181e+08 muA
** NormalTransistorNmos: 6.70124e+08 muA
** NormalTransistorPmos: -9.19049e+07 muA
** DiodeTransistorPmos: -5.33309e+07 muA
** NormalTransistorPmos: -5.33319e+07 muA
** NormalTransistorPmos: -5.33309e+07 muA
** DiodeTransistorPmos: -5.33319e+07 muA
** NormalTransistorNmos: 1.0666e+08 muA
** DiodeTransistorNmos: 1.06659e+08 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 1.17892e+09 muA
** NormalTransistorPmos: -1.17891e+09 muA
** NormalTransistorPmos: -1.17891e+09 muA
** DiodeTransistorNmos: 9.19041e+07 muA
** NormalTransistorNmos: 9.19041e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.9718e+08 muA
** DiodeTransistorPmos: -6.70123e+08 muA


** Expected Voltages: 
** ibias: 0.670001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.15901  V
** out: 2.5  V
** outFirstStage: 4.01601  V
** outInputVoltageBiasXXnXX1: 1.16201  V
** outSourceVoltageBiasXXnXX1: 0.581001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.27801  V
** innerTransistorStack1Load1: 4.27601  V
** out1: 3.46401  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.58001  V
** inner: 0.581001  V


.END