** Name: two_stage_single_output_op_amp_57_5

.MACRO two_stage_single_output_op_amp_57_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=5e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=126e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=4e-6 W=53e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=6e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=558e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=437e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=9e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=35e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=35e-6
mMainBias11 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=125e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=265e-6
mFoldedCascodeFirstStageLoad13 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=9e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=82e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=34e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=34e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=4e-6 W=153e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=6e-6
mSecondStage1StageBias20 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=558e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=126e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_57_5

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 5.65401 mW
** Area: 9772 (mu_m)^2
** Transit frequency: 4.16101 MHz
** Transit frequency with error factor: 4.15641 MHz
** Slew rate: 5.04532 V/mu_s
** Phase margin: 72.7657°
** CMRR: 103 dB
** VoutMax: 3.38001 V
** VoutMin: 0.570001 V
** VcmMax: 3.24001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 9.86401e+06 muA
** NormalTransistorNmos: 1.24238e+08 muA
** NormalTransistorNmos: 2.28241e+07 muA
** NormalTransistorNmos: 3.43351e+07 muA
** NormalTransistorNmos: 2.28241e+07 muA
** NormalTransistorNmos: 3.43351e+07 muA
** DiodeTransistorPmos: -2.28249e+07 muA
** NormalTransistorPmos: -2.28249e+07 muA
** NormalTransistorPmos: -2.30249e+07 muA
** NormalTransistorPmos: -2.30259e+07 muA
** NormalTransistorPmos: -1.15119e+07 muA
** NormalTransistorPmos: -1.15119e+07 muA
** NormalTransistorNmos: 9.17955e+08 muA
** NormalTransistorPmos: -9.17954e+08 muA
** DiodeTransistorPmos: -9.17955e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.86499e+06 muA
** NormalTransistorPmos: -9.86599e+06 muA
** DiodeTransistorPmos: -1.24237e+08 muA
** DiodeTransistorPmos: -1.24238e+08 muA


** Expected Voltages: 
** ibias: 1.18001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.89401  V
** out: 2.5  V
** outFirstStage: 0.975001  V
** outInputVoltageBiasXXpXX1: 2.81601  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 3.90801  V
** outSourceVoltageBiasXXpXX2: 4.18501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 3.64101  V
** out1: 4.26101  V
** sourceGCC1: 0.529001  V
** sourceGCC2: 0.529001  V
** sourceTransconductance: 3.25801  V
** inner: 3.90301  V


.END