** Name: two_stage_single_output_op_amp_82_12

.MACRO two_stage_single_output_op_amp_82_12 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=35e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=35e-6
mMainBias3 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=8e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=372e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=577e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=35e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=9e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=9e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=17e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mMainBias14 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mSecondStage1StageBias15 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=372e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=35e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=122e-6
mFoldedCascodeFirstStageLoad19 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=100e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=100e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=100e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=567e-6
mSecondStage1Transconductor23 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=308e-6
mFoldedCascodeFirstStageLoad24 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=100e-6
mMainBias25 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=38e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_82_12

** Expected Performance Values: 
** Gain: 178 dB
** Power consumption: 3.45601 mW
** Area: 14987 (mu_m)^2
** Transit frequency: 4.00601 MHz
** Transit frequency with error factor: 4.00645 MHz
** Slew rate: 3.77583 V/mu_s
** Phase margin: 63.0254°
** CMRR: 148 dB
** VoutMax: 4.29001 V
** VoutMin: 0.890001 V
** VcmMax: 5.02001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 1.35361e+07 muA
** NormalTransistorNmos: 1.49706e+08 muA
** NormalTransistorPmos: -9.95599e+06 muA
** NormalTransistorPmos: -1.71429e+07 muA
** NormalTransistorPmos: -2.57129e+07 muA
** NormalTransistorPmos: -1.71469e+07 muA
** NormalTransistorPmos: -2.57189e+07 muA
** DiodeTransistorNmos: 1.71441e+07 muA
** NormalTransistorNmos: 1.71451e+07 muA
** NormalTransistorNmos: 1.71461e+07 muA
** DiodeTransistorNmos: 1.71451e+07 muA
** NormalTransistorNmos: 1.71411e+07 muA
** DiodeTransistorNmos: 1.71401e+07 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 4.56478e+08 muA
** DiodeTransistorNmos: 4.56479e+08 muA
** NormalTransistorPmos: -4.56477e+08 muA
** NormalTransistorPmos: -4.56478e+08 muA
** DiodeTransistorNmos: 9.95701e+06 muA
** NormalTransistorNmos: 9.95801e+06 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.35369e+07 muA
** DiodeTransistorPmos: -1.49705e+08 muA


** Expected Voltages: 
** ibias: 1.29201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.22301  V
** outInputVoltageBiasXXnXX1: 1.24601  V
** outSourceVoltageBiasXXnXX1: 0.623001  V
** outSourceVoltageBiasXXnXX2: 0.647001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.05501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.633001  V
** innerTransistorStack2Load2: 0.633001  V
** out1: 1.19001  V
** sourceGCC1: 4.41901  V
** sourceGCC2: 4.41901  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.74701  V
** inner: 0.624001  V
** inner: 0.643001  V


.END