** Name: two_stage_single_output_op_amp_45_10

.MACRO two_stage_single_output_op_amp_45_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=46e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=119e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=54e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=59e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=59e-6
mSecondStage1StageBias9 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=597e-6
mFoldedCascodeFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=54e-6
mMainBias11 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=52e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=119e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=147e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=147e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=448e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
mMainBias17 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=449e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad19 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=84e-6
mMainBias20 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=424e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.2001e-12
.EOM two_stage_single_output_op_amp_45_10

** Expected Performance Values: 
** Gain: 135 dB
** Power consumption: 11.0131 mW
** Area: 8306 (mu_m)^2
** Transit frequency: 9.68001 MHz
** Transit frequency with error factor: 9.67982 MHz
** Slew rate: 6.52318 V/mu_s
** Phase margin: 60.1606°
** CMRR: 142 dB
** VoutMax: 4.25 V
** VoutMin: 0.170001 V
** VcmMax: 4.04001 V
** VcmMin: -0.389999 V


** Expected Currents: 
** NormalTransistorNmos: 1.31994e+08 muA
** NormalTransistorPmos: -1.21251e+08 muA
** NormalTransistorPmos: -1.15387e+08 muA
** NormalTransistorNmos: 8.63371e+07 muA
** NormalTransistorNmos: 1.48009e+08 muA
** NormalTransistorNmos: 8.63341e+07 muA
** NormalTransistorNmos: 1.48004e+08 muA
** DiodeTransistorPmos: -8.63359e+07 muA
** NormalTransistorPmos: -8.63349e+07 muA
** NormalTransistorPmos: -8.63359e+07 muA
** NormalTransistorPmos: -1.23338e+08 muA
** NormalTransistorPmos: -6.16699e+07 muA
** NormalTransistorPmos: -6.16699e+07 muA
** NormalTransistorNmos: 1.51794e+09 muA
** NormalTransistorPmos: -1.51793e+09 muA
** NormalTransistorPmos: -1.51793e+09 muA
** DiodeTransistorNmos: 1.21252e+08 muA
** DiodeTransistorNmos: 1.15388e+08 muA
** DiodeTransistorPmos: -1.31993e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.972001  V
** out: 2.5  V
** outFirstStage: 4.06101  V
** outVoltageBiasXXnXX2: 0.578001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.48901  V
** out1: 4.23401  V
** sourceGCC1: 0.373001  V
** sourceGCC2: 0.373001  V
** sourceTransconductance: 3.21701  V
** innerTransconductance: 4.625  V


.END