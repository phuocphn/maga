** Name: two_stage_single_output_op_amp_75_2

.MACRO two_stage_single_output_op_amp_75_2 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=25e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=543e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=25e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=11e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=536e-6
mSecondStage1Transconductor12 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=98e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=11e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=58e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=169e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=100e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=63e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=63e-6
mMainBias19 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=581e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=423e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=100e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_75_2

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 4.79601 mW
** Area: 14187 (mu_m)^2
** Transit frequency: 3.95101 MHz
** Transit frequency with error factor: 3.95139 MHz
** Slew rate: 4.70387 V/mu_s
** Phase margin: 63.0254°
** CMRR: 144 dB
** VoutMax: 4.62001 V
** VoutMin: 0.360001 V
** VcmMax: 5.03001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorNmos: 9.64561e+07 muA
** NormalTransistorNmos: 2.76506e+08 muA
** NormalTransistorPmos: -2.94724e+08 muA
** NormalTransistorPmos: -2.12689e+07 muA
** NormalTransistorPmos: -3.19019e+07 muA
** NormalTransistorPmos: -2.12719e+07 muA
** NormalTransistorPmos: -3.19069e+07 muA
** DiodeTransistorNmos: 2.12701e+07 muA
** NormalTransistorNmos: 2.12711e+07 muA
** NormalTransistorNmos: 2.12701e+07 muA
** NormalTransistorNmos: 2.12691e+07 muA
** NormalTransistorNmos: 2.12701e+07 muA
** NormalTransistorNmos: 1.06341e+07 muA
** NormalTransistorNmos: 1.06341e+07 muA
** NormalTransistorNmos: 2.17654e+08 muA
** NormalTransistorNmos: 2.17653e+08 muA
** NormalTransistorPmos: -2.17653e+08 muA
** DiodeTransistorNmos: 2.94725e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.64569e+07 muA
** DiodeTransistorPmos: -2.76505e+08 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.998001  V
** out: 2.5  V
** outFirstStage: 0.600001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.05801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.442001  V
** innerTransistorStack2Load2: 0.442001  V
** out1: 0.605001  V
** sourceGCC1: 4.40401  V
** sourceGCC2: 4.40401  V
** sourceTransconductance: 1.90501  V
** innerTransconductance: 0.431001  V


.END