** Name: two_stage_single_output_op_amp_79_8

.MACRO two_stage_single_output_op_amp_79_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=68e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=23e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=23e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=26e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=26e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=11e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=586e-6
mSecondStage1StageBias13 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=258e-6
mFoldedCascodeFirstStageLoad14 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=50e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=595e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=50e-6
mMainBias20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=504e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=87e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_79_8

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 7.13501 mW
** Area: 8001 (mu_m)^2
** Transit frequency: 4.16701 MHz
** Transit frequency with error factor: 4.16726 MHz
** Slew rate: 4.49538 V/mu_s
** Phase margin: 62.4525°
** CMRR: 140 dB
** VoutMax: 4.25 V
** VoutMin: 0.360001 V
** VcmMax: 5.17001 V
** VcmMin: 1.33001 V


** Expected Currents: 
** NormalTransistorPmos: -5.01631e+08 muA
** NormalTransistorPmos: -8.72709e+07 muA
** NormalTransistorPmos: -2.03059e+07 muA
** NormalTransistorPmos: -3.14299e+07 muA
** NormalTransistorPmos: -2.03059e+07 muA
** NormalTransistorPmos: -3.14299e+07 muA
** NormalTransistorNmos: 2.03051e+07 muA
** NormalTransistorNmos: 2.03041e+07 muA
** NormalTransistorNmos: 2.03051e+07 muA
** NormalTransistorNmos: 2.03041e+07 muA
** NormalTransistorNmos: 2.22451e+07 muA
** NormalTransistorNmos: 2.22441e+07 muA
** NormalTransistorNmos: 1.11231e+07 muA
** NormalTransistorNmos: 1.11231e+07 muA
** NormalTransistorNmos: 7.55159e+08 muA
** NormalTransistorNmos: 7.55158e+08 muA
** NormalTransistorPmos: -7.55158e+08 muA
** DiodeTransistorNmos: 5.01632e+08 muA
** DiodeTransistorNmos: 8.72701e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.10501  V
** outVoltageBiasXXnXX2: 0.580001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.545001  V
** innerTransistorStack1Load2: 0.545001  V
** innerTransistorStack2Load2: 0.545001  V
** out1: 0.727001  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.90601  V
** innerStageBias: 0.514001  V


.END