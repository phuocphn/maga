** Name: two_stage_single_output_op_amp_79_4

.MACRO two_stage_single_output_op_amp_79_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=213e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=85e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=103e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=103e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=33e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=71e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=71e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=25e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=91e-6
mSecondStage1Transconductor13 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=467e-6
mFoldedCascodeFirstStageLoad14 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=33e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=67e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=438e-6
mSecondStage1StageBias19 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=314e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=67e-6
mMainBias21 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=136e-6
mMainBias22 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=67e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.30001e-12
.EOM two_stage_single_output_op_amp_79_4

** Expected Performance Values: 
** Gain: 179 dB
** Power consumption: 3.74201 mW
** Area: 8362 (mu_m)^2
** Transit frequency: 5.38901 MHz
** Transit frequency with error factor: 5.38904 MHz
** Slew rate: 5.07669 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 3.92001 V
** VoutMin: 0.520001 V
** VcmMax: 5.17001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorPmos: -1.35948e+08 muA
** NormalTransistorPmos: -6.79289e+07 muA
** NormalTransistorPmos: -2.70329e+07 muA
** NormalTransistorPmos: -4.05549e+07 muA
** NormalTransistorPmos: -2.70329e+07 muA
** NormalTransistorPmos: -4.05549e+07 muA
** NormalTransistorNmos: 2.70321e+07 muA
** NormalTransistorNmos: 2.70311e+07 muA
** NormalTransistorNmos: 2.70321e+07 muA
** NormalTransistorNmos: 2.70311e+07 muA
** NormalTransistorNmos: 2.70451e+07 muA
** NormalTransistorNmos: 2.70441e+07 muA
** NormalTransistorNmos: 1.35231e+07 muA
** NormalTransistorNmos: 1.35231e+07 muA
** NormalTransistorNmos: 4.43431e+08 muA
** NormalTransistorNmos: 4.43432e+08 muA
** NormalTransistorPmos: -4.4343e+08 muA
** NormalTransistorPmos: -4.43431e+08 muA
** DiodeTransistorNmos: 1.35949e+08 muA
** DiodeTransistorNmos: 6.79281e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.746001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.951001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.350001  V
** innerTransistorStack1Load2: 0.375  V
** innerTransistorStack2Load2: 0.376001  V
** out1: 0.581001  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 4.25301  V
** innerTransconductance: 0.362001  V


.END