** Name: two_stage_single_output_op_amp_9_7

.MACRO two_stage_single_output_op_amp_9_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=22e-6
mSimpleFirstStageTransconductor3 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=8e-6
mSimpleFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mSecondStage1StageBias5 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=221e-6
mSimpleFirstStageTransconductor6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=8e-6
mSimpleFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=22e-6
mSecondStage1Transconductor8 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=38e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_9_7

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 2.38901 mW
** Area: 1181 (mu_m)^2
** Transit frequency: 2.86701 MHz
** Transit frequency with error factor: 2.86308 MHz
** Slew rate: 5.52777 V/mu_s
** Phase margin: 60.1606°
** CMRR: 101 dB
** negPSRR: 97 dB
** posPSRR: 88 dB
** VoutMax: 4.25 V
** VoutMin: 0.260001 V
** VcmMax: 4.21001 V
** VcmMin: 0.980001 V


** Expected Currents: 
** NormalTransistorPmos: -1.27529e+07 muA
** NormalTransistorPmos: -1.27529e+07 muA
** DiodeTransistorPmos: -1.27529e+07 muA
** NormalTransistorNmos: 2.55051e+07 muA
** NormalTransistorNmos: 1.27521e+07 muA
** NormalTransistorNmos: 1.27521e+07 muA
** NormalTransistorNmos: 4.42339e+08 muA
** NormalTransistorPmos: -4.42338e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA


** Expected Voltages: 
** ibias: 0.670001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.99501  V
** out1: 3.23801  V
** sourceTransconductance: 1.78701  V


.END