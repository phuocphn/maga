** Name: two_stage_single_output_op_amp_43_11

.MACRO two_stage_single_output_op_amp_43_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=12e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=172e-6
mSecondStage1StageBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=9e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=73e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=377e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=377e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=559e-6
mSecondStage1StageBias10 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=6e-6 W=126e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=73e-6
mMainBias12 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=94e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=370e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=427e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=449e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=172e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_43_11

** Expected Performance Values: 
** Gain: 133 dB
** Power consumption: 2.31601 mW
** Area: 13533 (mu_m)^2
** Transit frequency: 4.17901 MHz
** Transit frequency with error factor: 4.15685 MHz
** Slew rate: 7.33264 V/mu_s
** Phase margin: 60.7336°
** CMRR: 93 dB
** VoutMax: 4.70001 V
** VoutMin: 0.880001 V
** VcmMax: 3.52001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.05431e+07 muA
** NormalTransistorNmos: 1.94901e+06 muA
** NormalTransistorNmos: 7.99461e+07 muA
** NormalTransistorNmos: 1.20076e+08 muA
** NormalTransistorNmos: 7.99461e+07 muA
** NormalTransistorNmos: 1.20076e+08 muA
** DiodeTransistorPmos: -7.99469e+07 muA
** NormalTransistorPmos: -7.99469e+07 muA
** NormalTransistorPmos: -8.02609e+07 muA
** NormalTransistorPmos: -4.01299e+07 muA
** NormalTransistorPmos: -4.01299e+07 muA
** NormalTransistorNmos: 1.80532e+08 muA
** NormalTransistorNmos: 1.80531e+08 muA
** NormalTransistorPmos: -1.80531e+08 muA
** NormalTransistorPmos: -1.80532e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.05439e+07 muA
** DiodeTransistorPmos: -1.94999e+06 muA


** Expected Voltages: 
** ibias: 1.20301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.28201  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outVoltageBiasXXpXX1: 4.02101  V
** outVoltageBiasXXpXX2: 4.18901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.27401  V
** sourceGCC1: 0.518001  V
** sourceGCC2: 0.518001  V
** sourceTransconductance: 3.73101  V
** innerStageBias: 0.478001  V
** innerTransconductance: 4.73501  V


.END