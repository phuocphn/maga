** Name: two_stage_single_output_op_amp_77_9

.MACRO two_stage_single_output_op_amp_77_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=12e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=8e-6 W=9e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=37e-6
mMainBias4 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=10e-6 W=10e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=210e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=17e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=16e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=8e-6 W=9e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=18e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=37e-6
mSecondStage1StageBias15 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=210e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=12e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerOutputLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mMainBias20 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=129e-6
mMainBias21 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mSecondStage1Transconductor22 out outFirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=595e-6
mFoldedCascodeFirstStageLoad23 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=40e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_77_9

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 4.87801 mW
** Area: 10483 (mu_m)^2
** Transit frequency: 3.91401 MHz
** Transit frequency with error factor: 3.91378 MHz
** Slew rate: 3.59837 V/mu_s
** Phase margin: 64.1713°
** CMRR: 139 dB
** VoutMax: 4.25 V
** VoutMin: 1.64001 V
** VcmMax: 5.17001 V
** VcmMin: 1.69001 V


** Expected Currents: 
** NormalTransistorPmos: -1.30745e+08 muA
** NormalTransistorPmos: -1.90539e+07 muA
** NormalTransistorPmos: -1.62449e+07 muA
** NormalTransistorPmos: -2.53459e+07 muA
** NormalTransistorPmos: -1.62449e+07 muA
** NormalTransistorPmos: -2.53459e+07 muA
** DiodeTransistorNmos: 1.62441e+07 muA
** DiodeTransistorNmos: 1.62431e+07 muA
** NormalTransistorNmos: 1.62441e+07 muA
** NormalTransistorNmos: 1.62431e+07 muA
** NormalTransistorNmos: 1.81991e+07 muA
** NormalTransistorNmos: 1.81981e+07 muA
** NormalTransistorNmos: 9.10001e+06 muA
** NormalTransistorNmos: 9.10001e+06 muA
** NormalTransistorNmos: 7.55159e+08 muA
** DiodeTransistorNmos: 7.55158e+08 muA
** NormalTransistorPmos: -7.55158e+08 muA
** DiodeTransistorNmos: 1.30746e+08 muA
** NormalTransistorNmos: 1.30747e+08 muA
** DiodeTransistorNmos: 1.90531e+07 muA
** DiodeTransistorNmos: 1.90521e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.04201  V
** inputVoltageBiasXXnXX2: 1.64801  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 1.02101  V
** outSourceVoltageBiasXXnXX2: 0.770001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.57701  V
** innerStageBias: 0.896001  V
** innerTransistorStack1Load2: 0.816001  V
** innerTransistorStack2Load2: 0.813001  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.93101  V
** inner: 1.02201  V


.END