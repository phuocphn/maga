** Name: two_stage_single_output_op_amp_75_8

.MACRO two_stage_single_output_op_amp_75_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=77e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=19e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=26e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=77e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=27e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=27e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=39e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=589e-6
mSecondStage1StageBias12 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=543e-6
mFoldedCascodeFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=19e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=138e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=72e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=72e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=361e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=138e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=528e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=160e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_75_8

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 6.27501 mW
** Area: 11854 (mu_m)^2
** Transit frequency: 3.77801 MHz
** Transit frequency with error factor: 3.77817 MHz
** Slew rate: 4.0099 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 0.550001 V
** VcmMax: 5.15001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorPmos: -2.01467e+08 muA
** NormalTransistorPmos: -6.11909e+07 muA
** NormalTransistorPmos: -1.86329e+07 muA
** NormalTransistorPmos: -2.79489e+07 muA
** NormalTransistorPmos: -1.86329e+07 muA
** NormalTransistorPmos: -2.79489e+07 muA
** DiodeTransistorNmos: 1.86321e+07 muA
** NormalTransistorNmos: 1.86321e+07 muA
** NormalTransistorNmos: 1.86321e+07 muA
** NormalTransistorNmos: 1.86331e+07 muA
** NormalTransistorNmos: 1.86321e+07 muA
** NormalTransistorNmos: 9.31701e+06 muA
** NormalTransistorNmos: 9.31701e+06 muA
** NormalTransistorNmos: 9.16345e+08 muA
** NormalTransistorNmos: 9.16344e+08 muA
** NormalTransistorPmos: -9.16344e+08 muA
** DiodeTransistorNmos: 2.01468e+08 muA
** DiodeTransistorNmos: 6.11901e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.18201  V
** outVoltageBiasXXnXX1: 1.15401  V
** outVoltageBiasXXnXX2: 0.639001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.581001  V
** innerTransistorStack2Load2: 0.508001  V
** out1: 0.574001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.92601  V
** innerStageBias: 0.434001  V


.END