** Name: two_stage_single_output_op_amp_12_12

.MACRO two_stage_single_output_op_amp_12_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=9e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=279e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=55e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=284e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=120e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=9e-6
mSecondStage1StageBias9 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=279e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=284e-6
mMainBias11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=31e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=101e-6
mSimpleFirstStageLoad13 FirstStageYinnerSourceLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=99e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=22e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=22e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=583e-6
mSecondStage1Transconductor17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad18 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=99e-6
mMainBias19 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=84e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.9001e-12
.EOM two_stage_single_output_op_amp_12_12

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 9.04601 mW
** Area: 10396 (mu_m)^2
** Transit frequency: 11.5981 MHz
** Transit frequency with error factor: 11.5918 MHz
** Slew rate: 10.9306 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** negPSRR: 108 dB
** posPSRR: 100 dB
** VoutMax: 4.25 V
** VoutMin: 1.53001 V
** VcmMax: 4.85001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorNmos: 3.12281e+07 muA
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -4.74809e+07 muA
** NormalTransistorPmos: -6.01029e+07 muA
** NormalTransistorPmos: -6.01039e+07 muA
** NormalTransistorPmos: -6.01029e+07 muA
** NormalTransistorPmos: -6.01039e+07 muA
** NormalTransistorNmos: 1.20204e+08 muA
** NormalTransistorNmos: 6.01021e+07 muA
** NormalTransistorNmos: 6.01021e+07 muA
** NormalTransistorNmos: 1.49874e+09 muA
** DiodeTransistorNmos: 1.49874e+09 muA
** NormalTransistorPmos: -1.49873e+09 muA
** NormalTransistorPmos: -1.49874e+09 muA
** DiodeTransistorNmos: 4.74801e+07 muA
** NormalTransistorNmos: 4.74801e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.12289e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 0.593001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.05801  V
** outInputVoltageBiasXXnXX1: 1.93201  V
** outSourceVoltageBiasXXnXX1: 0.966001  V
** outVoltageBiasXXpXX0: 4.25801  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.88201  V
** innerTransistorStack1Load1: 4.43401  V
** innerTransistorStack2Load1: 4.43401  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.62201  V
** inner: 0.966001  V


.END