** Name: two_stage_single_output_op_amp_82_10

.MACRO two_stage_single_output_op_amp_82_10 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=3e-6 W=85e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=85e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=39e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=215e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=3e-6 W=85e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=56e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=56e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=39e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias13 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=599e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=85e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=93e-6
mMainBias16 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=36e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=241e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=466e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=466e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=388e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=591e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=241e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=110e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.7001e-12
.EOM two_stage_single_output_op_amp_82_10

** Expected Performance Values: 
** Gain: 134 dB
** Power consumption: 8.99101 mW
** Area: 10617 (mu_m)^2
** Transit frequency: 5.44301 MHz
** Transit frequency with error factor: 5.44327 MHz
** Slew rate: 4.70782 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 4.25 V
** VoutMin: 0.310001 V
** VcmMax: 5.14001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorNmos: 1.82761e+08 muA
** NormalTransistorNmos: 7.06311e+07 muA
** NormalTransistorPmos: -3.56169e+07 muA
** NormalTransistorPmos: -9.78779e+07 muA
** NormalTransistorPmos: -1.51208e+08 muA
** NormalTransistorPmos: -9.78779e+07 muA
** NormalTransistorPmos: -1.51208e+08 muA
** DiodeTransistorNmos: 9.78771e+07 muA
** NormalTransistorNmos: 9.78761e+07 muA
** NormalTransistorNmos: 9.78771e+07 muA
** DiodeTransistorNmos: 9.78761e+07 muA
** NormalTransistorNmos: 1.0666e+08 muA
** DiodeTransistorNmos: 1.06659e+08 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 1.19687e+09 muA
** NormalTransistorPmos: -1.19686e+09 muA
** NormalTransistorPmos: -1.19686e+09 muA
** DiodeTransistorNmos: 3.56161e+07 muA
** NormalTransistorNmos: 3.56151e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.8276e+08 muA
** DiodeTransistorPmos: -7.06319e+07 muA


** Expected Voltages: 
** ibias: 0.711001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.02101  V
** outInputVoltageBiasXXnXX1: 1.16801  V
** outSourceVoltageBiasXXnXX1: 0.584001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.16601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.606001  V
** innerTransistorStack2Load2: 0.606001  V
** out1: 1.17601  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.58501  V
** inner: 0.583001  V


.END