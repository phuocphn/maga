** Name: two_stage_single_output_op_amp_44_11

.MACRO two_stage_single_output_op_amp_44_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=8e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=387e-6
mSecondStage1StageBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=11e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=29e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=107e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=107e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSecondStage1StageBias10 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=260e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=29e-6
mMainBias12 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=155e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=387e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=96e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=96e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=78e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=508e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=597e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=224e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.80001e-12
.EOM two_stage_single_output_op_amp_44_11

** Expected Performance Values: 
** Gain: 167 dB
** Power consumption: 3.29201 mW
** Area: 13613 (mu_m)^2
** Transit frequency: 3.45401 MHz
** Transit frequency with error factor: 3.45438 MHz
** Slew rate: 7.87685 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 4.29001 V
** VoutMin: 0.790001 V
** VcmMax: 3.61001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorNmos: 6.67101e+06 muA
** NormalTransistorNmos: 4.62791e+07 muA
** NormalTransistorNmos: 6.99771e+07 muA
** NormalTransistorNmos: 4.62791e+07 muA
** NormalTransistorNmos: 6.99771e+07 muA
** NormalTransistorPmos: -4.62799e+07 muA
** NormalTransistorPmos: -4.62799e+07 muA
** DiodeTransistorPmos: -4.62799e+07 muA
** NormalTransistorPmos: -4.73989e+07 muA
** NormalTransistorPmos: -2.36989e+07 muA
** NormalTransistorPmos: -2.36989e+07 muA
** NormalTransistorNmos: 4.00319e+08 muA
** NormalTransistorNmos: 4.00318e+08 muA
** NormalTransistorPmos: -4.00318e+08 muA
** NormalTransistorPmos: -4.00319e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -6.67199e+06 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.92001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 3.98301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.27201  V
** out1: 3.55601  V
** sourceGCC1: 0.529001  V
** sourceGCC2: 0.529001  V
** sourceTransconductance: 3.43401  V
** innerStageBias: 0.534001  V
** innerTransconductance: 4.44301  V


.END