** Name: two_stage_single_output_op_amp_48_10

.MACRO two_stage_single_output_op_amp_48_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=88e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=481e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=481e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=314e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=193e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=193e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=555e-6
mFoldedCascodeFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=314e-6
mMainBias12 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=190e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=481e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=22e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=22e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=548e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=105e-6
mMainBias18 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=112e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=481e-6
mMainBias21 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=306e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.6001e-12
.EOM two_stage_single_output_op_amp_48_10

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 6.06801 mW
** Area: 14969 (mu_m)^2
** Transit frequency: 2.66301 MHz
** Transit frequency with error factor: 2.66278 MHz
** Slew rate: 9.2599 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 4.25 V
** VoutMin: 0.150001 V
** VcmMax: 3.44001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.82761e+08 muA
** NormalTransistorPmos: -3.08339e+07 muA
** NormalTransistorPmos: -8.38049e+07 muA
** NormalTransistorNmos: 1.09341e+08 muA
** NormalTransistorNmos: 1.83798e+08 muA
** NormalTransistorNmos: 1.09341e+08 muA
** NormalTransistorNmos: 1.83798e+08 muA
** DiodeTransistorPmos: -1.0934e+08 muA
** NormalTransistorPmos: -1.09341e+08 muA
** NormalTransistorPmos: -1.0934e+08 muA
** DiodeTransistorPmos: -1.09341e+08 muA
** NormalTransistorPmos: -1.48916e+08 muA
** NormalTransistorPmos: -7.44579e+07 muA
** NormalTransistorPmos: -7.44579e+07 muA
** NormalTransistorNmos: 5.28535e+08 muA
** NormalTransistorPmos: -5.28534e+08 muA
** NormalTransistorPmos: -5.28535e+08 muA
** DiodeTransistorNmos: 3.08331e+07 muA
** DiodeTransistorNmos: 8.38041e+07 muA
** DiodeTransistorPmos: -1.8276e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.926001  V
** out: 2.5  V
** outFirstStage: 3.90701  V
** outVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.27601  V
** innerTransistorStack1Load2: 4.27501  V
** out1: 3.55201  V
** sourceGCC1: 0.364001  V
** sourceGCC2: 0.364001  V
** sourceTransconductance: 3.81401  V
** innerTransconductance: 4.47101  V


.END