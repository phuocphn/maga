** Name: two_stage_single_output_op_amp_15_1

.MACRO two_stage_single_output_op_amp_15_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=33e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=46e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=63e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=21e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=198e-6
mSimpleFirstStageLoad7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=33e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=157e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=12e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=21e-6
mMainBias11 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=550e-6
mSecondStage1StageBias12 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=585e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=12e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_15_1

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 1.33701 mW
** Area: 5334 (mu_m)^2
** Transit frequency: 2.58901 MHz
** Transit frequency with error factor: 2.58133 MHz
** Slew rate: 3.83957 V/mu_s
** Phase margin: 64.1713°
** CMRR: 94 dB
** negPSRR: 96 dB
** posPSRR: 148 dB
** VoutMax: 4.84001 V
** VoutMin: 0.150001 V
** VcmMax: 3.11001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 3.99981e+07 muA
** NormalTransistorPmos: -8.76139e+07 muA
** DiodeTransistorNmos: 1.25711e+07 muA
** NormalTransistorNmos: 1.25711e+07 muA
** NormalTransistorPmos: -2.51449e+07 muA
** NormalTransistorPmos: -2.51459e+07 muA
** NormalTransistorPmos: -1.25719e+07 muA
** NormalTransistorPmos: -1.25719e+07 muA
** NormalTransistorNmos: 9.46681e+07 muA
** NormalTransistorPmos: -9.46689e+07 muA
** DiodeTransistorNmos: 8.76131e+07 muA
** DiodeTransistorPmos: -3.99989e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.555001  V
** inputVoltageBiasXXpXX1: 3.98301  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.80501  V
** out1: 0.555001  V
** sourceTransconductance: 3.40501  V


.END