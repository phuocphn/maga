** Name: two_stage_single_output_op_amp_148_9

.MACRO two_stage_single_output_op_amp_148_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=45e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=3e-6 W=23e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=5e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=186e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=32e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=14e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=3e-6 W=23e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=50e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=186e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=45e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=14e-6
mSimpleFirstStageLoad15 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=202e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=366e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=366e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=411e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=202e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_148_9

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 7.36701 mW
** Area: 6875 (mu_m)^2
** Transit frequency: 2.76801 MHz
** Transit frequency with error factor: 2.76557 MHz
** Slew rate: 3.50015 V/mu_s
** Phase margin: 69.9009°
** CMRR: 126 dB
** VoutMax: 4.25 V
** VoutMin: 1.33001 V
** VcmMax: 4.85001 V
** VcmMin: 0.790001 V


** Expected Currents: 
** NormalTransistorPmos: -1.82489e+07 muA
** NormalTransistorPmos: -1.01379e+07 muA
** DiodeTransistorNmos: 3.61184e+08 muA
** DiodeTransistorNmos: 3.61183e+08 muA
** NormalTransistorNmos: 3.61182e+08 muA
** NormalTransistorNmos: 3.61183e+08 muA
** NormalTransistorPmos: -3.69182e+08 muA
** NormalTransistorPmos: -3.69181e+08 muA
** NormalTransistorPmos: -3.6918e+08 muA
** NormalTransistorPmos: -3.69181e+08 muA
** NormalTransistorNmos: 1.59991e+07 muA
** NormalTransistorNmos: 7.99901e+06 muA
** NormalTransistorNmos: 7.99901e+06 muA
** NormalTransistorNmos: 6.86587e+08 muA
** DiodeTransistorNmos: 6.86586e+08 muA
** NormalTransistorPmos: -6.86586e+08 muA
** DiodeTransistorNmos: 1.82481e+07 muA
** NormalTransistorNmos: 1.82471e+07 muA
** DiodeTransistorNmos: 1.01371e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.74001  V
** outSourceVoltageBiasXXnXX1: 0.870001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.589001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerTransistorStack1Load1: 1.15401  V
** innerTransistorStack1Load2: 4.29201  V
** innerTransistorStack2Load1: 1.15501  V
** innerTransistorStack2Load2: 4.29201  V
** sourceTransconductance: 1.89301  V
** inner: 0.869001  V


.END