** Name: two_stage_single_output_op_amp_170_3

.MACRO two_stage_single_output_op_amp_170_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=49e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=8e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=8e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=35e-6
mMainBias6 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=8e-6 W=8e-6
mSimpleFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=125e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
mSimpleFirstStageLoad9 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=10e-6 W=148e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=148e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=148e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=150e-6
mSimpleFirstStageLoad13 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=148e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=35e-6
mMainBias15 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=53e-6
mSimpleFirstStageTransconductor16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=15e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=8e-6
mSimpleFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=125e-6
mSecondStage1StageBias19 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=231e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=35e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=8e-6 W=296e-6
mSimpleFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=5e-6 W=8e-6
mSimpleFirstStageTransconductor23 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=15e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.40001e-12
.EOM two_stage_single_output_op_amp_170_3

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 1.87801 mW
** Area: 14864 (mu_m)^2
** Transit frequency: 2.78201 MHz
** Transit frequency with error factor: 2.78019 MHz
** Slew rate: 3.69049 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 3.02001 V
** VoutMin: 0.300001 V
** VcmMax: 3.15001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 6.66701e+06 muA
** NormalTransistorNmos: 1.01511e+07 muA
** DiodeTransistorPmos: -1.62449e+07 muA
** DiodeTransistorPmos: -1.62449e+07 muA
** NormalTransistorPmos: -1.62449e+07 muA
** NormalTransistorPmos: -1.62449e+07 muA
** NormalTransistorNmos: 2.81891e+07 muA
** NormalTransistorNmos: 2.81891e+07 muA
** NormalTransistorNmos: 2.81891e+07 muA
** NormalTransistorNmos: 2.81891e+07 muA
** NormalTransistorPmos: -2.38909e+07 muA
** DiodeTransistorPmos: -2.38919e+07 muA
** NormalTransistorPmos: -1.19449e+07 muA
** NormalTransistorPmos: -1.19449e+07 muA
** NormalTransistorNmos: 2.92374e+08 muA
** NormalTransistorPmos: -2.92373e+08 muA
** NormalTransistorPmos: -2.92374e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -6.66799e+06 muA
** NormalTransistorPmos: -6.66899e+06 muA
** DiodeTransistorPmos: -1.01519e+07 muA
** DiodeTransistorPmos: -1.01529e+07 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.710001  V
** outInputVoltageBiasXXpXX1: 3.36401  V
** outInputVoltageBiasXXpXX2: 2.37201  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.18201  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerSourceLoad1: 3.68601  V
** innerTransistorStack1Load2: 0.560001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.560001  V
** sourceTransconductance: 3.27501  V
** innerStageBias: 3.59801  V
** inner: 4.18001  V


.END