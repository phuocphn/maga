** Name: one_stage_single_output_op_amp67

.MACRO one_stage_single_output_op_amp67 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=317e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=249e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=7e-6 W=225e-6
mFoldedCascodeFirstStageLoad4 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=225e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=21e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerOutputLoad2 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=159e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=188e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=188e-6
mFoldedCascodeFirstStageLoad10 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=159e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=308e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=225e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=387e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=387e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=327e-6
mMainBias16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad17 out FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=225e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp67

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 7.70901 mW
** Area: 7350 (mu_m)^2
** Transit frequency: 16.4651 MHz
** Transit frequency with error factor: 16.4646 MHz
** Slew rate: 15.0743 V/mu_s
** Phase margin: 88.8085°
** CMRR: 129 dB
** VoutMax: 3.32001 V
** VoutMin: 0.720001 V
** VcmMax: 3.25 V
** VcmMin: -0.389999 V


** Expected Currents: 
** NormalTransistorPmos: -6.03767e+08 muA
** NormalTransistorNmos: 3.02837e+08 muA
** NormalTransistorNmos: 4.58973e+08 muA
** NormalTransistorNmos: 3.02837e+08 muA
** NormalTransistorNmos: 4.58973e+08 muA
** DiodeTransistorPmos: -3.02836e+08 muA
** NormalTransistorPmos: -3.02837e+08 muA
** NormalTransistorPmos: -3.02836e+08 muA
** DiodeTransistorPmos: -3.02837e+08 muA
** NormalTransistorPmos: -3.12274e+08 muA
** NormalTransistorPmos: -3.12273e+08 muA
** NormalTransistorPmos: -1.56136e+08 muA
** NormalTransistorPmos: -1.56136e+08 muA
** DiodeTransistorNmos: 6.03768e+08 muA
** DiodeTransistorNmos: 6.03767e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.12901  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.574001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 2.75301  V
** innerStageBias: 4.26601  V
** innerTransistorStack1Load2: 4.04001  V
** innerTransistorStack2Load2: 4.04601  V
** sourceGCC1: 0.574001  V
** sourceGCC2: 0.574001  V
** sourceTransconductance: 3.21401  V


.END