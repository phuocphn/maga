** Name: two_stage_single_output_op_amp_76_12

.MACRO two_stage_single_output_op_amp_76_12 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=142e-6
mMainBias2 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=70e-6
mMainBias4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=6e-6 W=126e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=61e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=517e-6
mMainBias7 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mMainBias8 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mMainBias9 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=142e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=90e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=90e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=61e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=70e-6
mMainBias15 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=126e-6
mSecondStage1StageBias16 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=517e-6
mFoldedCascodeFirstStageLoad17 outFirstStage inputVoltageBiasXXnXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=36e-6
mMainBias18 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mFoldedCascodeFirstStageLoad19 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=178e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=273e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=273e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=481e-6
mMainBias23 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=155e-6
mSecondStage1Transconductor24 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad25 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=178e-6
mMainBias26 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=217e-6
mMainBias27 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=553e-6
mMainBias28 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=75e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.6001e-12
.EOM two_stage_single_output_op_amp_76_12

** Expected Performance Values: 
** Gain: 171 dB
** Power consumption: 11.9781 mW
** Area: 14987 (mu_m)^2
** Transit frequency: 7.27701 MHz
** Transit frequency with error factor: 7.27744 MHz
** Slew rate: 6.36746 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 1.26001 V
** VcmMax: 5.22001 V
** VcmMin: 1.90001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -4.43259e+07 muA
** NormalTransistorPmos: -1.29049e+08 muA
** NormalTransistorPmos: -3.25433e+08 muA
** NormalTransistorPmos: -9.14959e+07 muA
** NormalTransistorPmos: -1.06089e+08 muA
** NormalTransistorPmos: -1.63227e+08 muA
** NormalTransistorPmos: -1.06089e+08 muA
** NormalTransistorPmos: -1.63227e+08 muA
** DiodeTransistorNmos: 1.0609e+08 muA
** NormalTransistorNmos: 1.0609e+08 muA
** NormalTransistorNmos: 1.0609e+08 muA
** NormalTransistorNmos: 1.14278e+08 muA
** DiodeTransistorNmos: 1.14277e+08 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 1.35721e+09 muA
** DiodeTransistorNmos: 1.35721e+09 muA
** NormalTransistorPmos: -1.3572e+09 muA
** NormalTransistorPmos: -1.35721e+09 muA
** DiodeTransistorNmos: 4.43251e+07 muA
** DiodeTransistorNmos: 1.2905e+08 muA
** NormalTransistorNmos: 1.29049e+08 muA
** DiodeTransistorNmos: 3.25434e+08 muA
** NormalTransistorNmos: 3.25435e+08 muA
** DiodeTransistorNmos: 9.14951e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX3: 1.08901  V
** out: 2.5  V
** outFirstStage: 4.04001  V
** outInputVoltageBiasXXnXX1: 1.74801  V
** outInputVoltageBiasXXnXX2: 1.67001  V
** outSourceVoltageBiasXXnXX1: 0.874001  V
** outSourceVoltageBiasXXnXX2: 0.835001  V
** outVoltageBiasXXnXX0: 1.125  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.362001  V
** out1: 0.567001  V
** sourceGCC1: 4.43201  V
** sourceGCC2: 4.43201  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.60401  V
** inner: 0.874001  V
** inner: 0.836001  V


.END