** Name: two_stage_single_output_op_amp_117_8

.MACRO two_stage_single_output_op_amp_117_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=10e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=25e-6
mMainBias3 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mTelescopicFirstStageLoad4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=154e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=41e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=28e-6
mTelescopicFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=156e-6
mTelescopicFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=32e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=16e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=16e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=301e-6
mTelescopicFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=32e-6
mMainBias14 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=15e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=67e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=125e-6
mTelescopicFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=154e-6
mMainBias18 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=264e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=572e-6
mTelescopicFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=96e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.30001e-12
.EOM two_stage_single_output_op_amp_117_8

** Expected Performance Values: 
** Gain: 147 dB
** Power consumption: 4.23201 mW
** Area: 6428 (mu_m)^2
** Transit frequency: 8.81301 MHz
** Transit frequency with error factor: 8.81281 MHz
** Slew rate: 21.1553 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 4.76001 V
** VoutMin: 0.780001 V
** VcmMax: 4.14001 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorNmos: 1.48001e+07 muA
** NormalTransistorNmos: 6.58291e+07 muA
** NormalTransistorPmos: -9.42899e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** DiodeTransistorPmos: -3.04759e+07 muA
** NormalTransistorPmos: -3.04759e+07 muA
** NormalTransistorPmos: -3.04759e+07 muA
** NormalTransistorNmos: 1.55239e+08 muA
** NormalTransistorNmos: 1.55238e+08 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 6.00478e+08 muA
** NormalTransistorNmos: 6.00477e+08 muA
** NormalTransistorPmos: -6.00477e+08 muA
** DiodeTransistorNmos: 9.42891e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.48009e+07 muA
** DiodeTransistorPmos: -6.58299e+07 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.65001  V
** out: 2.5  V
** outFirstStage: 4.19301  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX0: 4.23601  V
** outVoltageBiasXXpXX1: 3.62901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.539001  V
** innerTransistorStack2Load2: 4.49001  V
** out1: 4.17701  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.493001  V


.END