** Name: two_stage_single_output_op_amp_121_12

.MACRO two_stage_single_output_op_amp_121_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=6e-6 W=26e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=160e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=562e-6
mMainBias4 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=10e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mTelescopicFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=158e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=34e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=17e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=17e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=160e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=562e-6
mTelescopicFirstStageLoad14 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=34e-6
mMainBias15 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=75e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=214e-6
mTelescopicFirstStageStageBias17 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=67e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=20e-6
mTelescopicFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=20e-6
mTelescopicFirstStageLoad20 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=14e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=474e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=599e-6
mTelescopicFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=14e-6
mMainBias24 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=211e-6
mMainBias25 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=13e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.30001e-12
.EOM two_stage_single_output_op_amp_121_12

** Expected Performance Values: 
** Gain: 177 dB
** Power consumption: 7.65801 mW
** Area: 9766 (mu_m)^2
** Transit frequency: 3.68901 MHz
** Transit frequency with error factor: 3.68892 MHz
** Slew rate: 5.50158 V/mu_s
** Phase margin: 62.4525°
** CMRR: 135 dB
** VoutMax: 3.76001 V
** VoutMin: 0.700001 V
** VcmMax: 4.58001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 2.42761e+07 muA
** NormalTransistorNmos: 6.93851e+07 muA
** NormalTransistorPmos: -3.06216e+08 muA
** NormalTransistorPmos: -1.88589e+07 muA
** NormalTransistorNmos: 1.61901e+07 muA
** NormalTransistorNmos: 1.61901e+07 muA
** NormalTransistorPmos: -1.61909e+07 muA
** NormalTransistorPmos: -1.61919e+07 muA
** NormalTransistorPmos: -1.61909e+07 muA
** NormalTransistorPmos: -1.61919e+07 muA
** NormalTransistorNmos: 5.12371e+07 muA
** NormalTransistorNmos: 5.12361e+07 muA
** NormalTransistorNmos: 1.61901e+07 muA
** NormalTransistorNmos: 1.61901e+07 muA
** NormalTransistorNmos: 1.07041e+09 muA
** DiodeTransistorNmos: 1.07041e+09 muA
** NormalTransistorPmos: -1.0704e+09 muA
** NormalTransistorPmos: -1.0704e+09 muA
** DiodeTransistorNmos: 3.06217e+08 muA
** NormalTransistorNmos: 3.06216e+08 muA
** DiodeTransistorNmos: 1.88581e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.42769e+07 muA
** DiodeTransistorPmos: -6.93859e+07 muA


** Expected Voltages: 
** ibias: 1.12601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.64101  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX3: 0.556001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 4.03501  V
** outVoltageBiasXXpXX1: 3.19601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.488001  V
** innerTransistorStack1Load2: 4.11801  V
** innerTransistorStack2Load2: 4.11801  V
** out1: 3.76001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.20501  V
** inner: 0.554001  V


.END