** Name: two_stage_single_output_op_amp_161_6

.MACRO two_stage_single_output_op_amp_161_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=17e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=65e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=1e-6 W=97e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=58e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=299e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=344e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=344e-6
mSimpleFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=346e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=589e-6
mMainBias12 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=115e-6
mSecondStage1Transconductor13 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=591e-6
mSimpleFirstStageLoad14 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=346e-6
mSimpleFirstStageStageBias15 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=369e-6
mSimpleFirstStageTransconductor16 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=248e-6
mSimpleFirstStageLoad17 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=1e-6 W=97e-6
mSimpleFirstStageStageBias18 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=185e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=58e-6
mSecondStage1StageBias20 out inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=299e-6
mSimpleFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=245e-6
mSimpleFirstStageTransconductor22 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=248e-6
mMainBias23 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=129e-6
mMainBias24 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=123e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14e-12
.EOM two_stage_single_output_op_amp_161_6

** Expected Performance Values: 
** Gain: 140 dB
** Power consumption: 14.6861 mW
** Area: 6687 (mu_m)^2
** Transit frequency: 14.4061 MHz
** Transit frequency with error factor: 14.3931 MHz
** Slew rate: 26.2989 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** VoutMax: 3.13001 V
** VoutMin: 0.300001 V
** VcmMax: 3.01001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 2.19033e+08 muA
** NormalTransistorPmos: -1.30789e+08 muA
** NormalTransistorPmos: -1.23801e+08 muA
** NormalTransistorPmos: -4.7194e+08 muA
** NormalTransistorPmos: -4.7194e+08 muA
** DiodeTransistorPmos: -4.7194e+08 muA
** NormalTransistorNmos: 6.59002e+08 muA
** NormalTransistorNmos: 6.59001e+08 muA
** NormalTransistorNmos: 6.59002e+08 muA
** NormalTransistorNmos: 6.59001e+08 muA
** NormalTransistorPmos: -3.74121e+08 muA
** NormalTransistorPmos: -3.7412e+08 muA
** NormalTransistorPmos: -1.8706e+08 muA
** NormalTransistorPmos: -1.8706e+08 muA
** NormalTransistorNmos: 1.12564e+09 muA
** NormalTransistorNmos: 1.12564e+09 muA
** NormalTransistorPmos: -1.12563e+09 muA
** DiodeTransistorPmos: -1.12563e+09 muA
** DiodeTransistorNmos: 1.3079e+08 muA
** DiodeTransistorNmos: 1.23802e+08 muA
** DiodeTransistorPmos: -2.19032e+08 muA
** NormalTransistorPmos: -2.19033e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 2.56801  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.78401  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX1: 0.705001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.29701  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load1: 3.91201  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 2.88201  V
** sourceTransconductance: 3.35401  V
** innerTransconductance: 0.150001  V
** inner: 3.77901  V


.END