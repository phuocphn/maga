** Name: two_stage_single_output_op_amp_74_7

.MACRO two_stage_single_output_op_amp_74_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=67e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=13e-6
mFoldedCascodeFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=34e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=18e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=10e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=24e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=67e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=10e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=34e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mSecondStage1StageBias12 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=191e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=8e-6 W=102e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=226e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=183e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=183e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=363e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=226e-6
mMainBias19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=58e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=139e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6e-12
.EOM two_stage_single_output_op_amp_74_7

** Expected Performance Values: 
** Gain: 112 dB
** Power consumption: 4.36701 mW
** Area: 7493 (mu_m)^2
** Transit frequency: 3.03501 MHz
** Transit frequency with error factor: 3.03525 MHz
** Slew rate: 7.53494 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 4.25 V
** VoutMin: 0.520001 V
** VcmMax: 5.19001 V
** VcmMin: 1.95001 V


** Expected Currents: 
** NormalTransistorPmos: -2.45139e+07 muA
** NormalTransistorPmos: -5.89969e+07 muA
** NormalTransistorPmos: -4.58929e+07 muA
** NormalTransistorPmos: -7.77729e+07 muA
** NormalTransistorPmos: -4.58929e+07 muA
** NormalTransistorPmos: -7.77729e+07 muA
** NormalTransistorNmos: 4.58921e+07 muA
** NormalTransistorNmos: 4.58921e+07 muA
** DiodeTransistorNmos: 4.58921e+07 muA
** NormalTransistorNmos: 6.37571e+07 muA
** DiodeTransistorNmos: 6.37561e+07 muA
** NormalTransistorNmos: 3.18791e+07 muA
** NormalTransistorNmos: 3.18791e+07 muA
** NormalTransistorNmos: 6.14281e+08 muA
** NormalTransistorPmos: -6.1428e+08 muA
** DiodeTransistorNmos: 2.45131e+07 muA
** NormalTransistorNmos: 2.45121e+07 muA
** DiodeTransistorNmos: 5.89961e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.40401  V
** outSourceVoltageBiasXXnXX1: 0.702001  V
** outSourceVoltageBiasXXpXX1: 4.21901  V
** outVoltageBiasXXnXX2: 0.923001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.561001  V
** out1: 1.17201  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.54401  V
** inner: 0.700001  V


.END