** Name: two_stage_single_output_op_amp_190_8

.MACRO two_stage_single_output_op_amp_190_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=8e-6 W=22e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=31e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=15e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=64e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=36e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=9e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=38e-6
mSimpleFirstStageLoad9 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=8e-6 W=22e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=16e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=174e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=31e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=252e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=33e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=38e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=126e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=126e-6
mSimpleFirstStageLoad18 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=253e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=377e-6
mSimpleFirstStageLoad20 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=253e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=28e-6
mMainBias22 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=307e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_190_8

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 8.17101 mW
** Area: 8081 (mu_m)^2
** Transit frequency: 3.71301 MHz
** Transit frequency with error factor: 3.7116 MHz
** Slew rate: 3.5001 V/mu_s
** Phase margin: 68.182°
** CMRR: 121 dB
** VoutMax: 4.25 V
** VoutMin: 0.870001 V
** VcmMax: 4.55001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorPmos: -3.12299e+07 muA
** NormalTransistorPmos: -3.46063e+08 muA
** NormalTransistorNmos: 1.3194e+08 muA
** NormalTransistorNmos: 1.31941e+08 muA
** DiodeTransistorNmos: 1.3194e+08 muA
** NormalTransistorPmos: -1.39981e+08 muA
** NormalTransistorPmos: -1.39982e+08 muA
** NormalTransistorPmos: -1.39982e+08 muA
** NormalTransistorPmos: -1.39982e+08 muA
** NormalTransistorNmos: 1.60851e+07 muA
** DiodeTransistorNmos: 1.60841e+07 muA
** NormalTransistorNmos: 8.04201e+06 muA
** NormalTransistorNmos: 8.04201e+06 muA
** NormalTransistorNmos: 9.56958e+08 muA
** NormalTransistorNmos: 9.56957e+08 muA
** NormalTransistorPmos: -9.56957e+08 muA
** DiodeTransistorNmos: 3.12291e+07 muA
** NormalTransistorNmos: 3.12281e+07 muA
** DiodeTransistorNmos: 3.46064e+08 muA
** DiodeTransistorNmos: 3.46063e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.12201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.18601  V
** outInputVoltageBiasXXnXX2: 1.58401  V
** outSourceVoltageBiasXXnXX1: 0.593001  V
** outSourceVoltageBiasXXnXX2: 0.659001  V
** outSourceVoltageBiasXXpXX1: 3.93501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.03701  V
** innerTransistorStack2Load1: 1.15501  V
** innerTransistorStack2Load2: 4.03701  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.967001  V
** inner: 0.592001  V


.END