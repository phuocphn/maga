** Name: two_stage_single_output_op_amp_97_7

.MACRO two_stage_single_output_op_amp_97_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=49e-6
mTelescopicFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=67e-6
mTelescopicFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=67e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=244e-6
mTelescopicFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=90e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=15e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=15e-6
mMainBias9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=314e-6
mSecondStage1StageBias10 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=90e-6
mTelescopicFirstStageStageBias12 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=122e-6
mTelescopicFirstStageLoad13 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=67e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=339e-6
mTelescopicFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=67e-6
mMainBias16 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20e-12
.EOM two_stage_single_output_op_amp_97_7

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 5.20701 mW
** Area: 4691 (mu_m)^2
** Transit frequency: 3.02501 MHz
** Transit frequency with error factor: 3.02469 MHz
** Slew rate: 5.97089 V/mu_s
** Phase margin: 60.1606°
** CMRR: 150 dB
** VoutMax: 4.68001 V
** VoutMin: 0.150001 V
** VcmMax: 3.82001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorNmos: 3.11332e+08 muA
** NormalTransistorPmos: -6.25399e+07 muA
** NormalTransistorNmos: 2.85711e+07 muA
** NormalTransistorNmos: 2.85711e+07 muA
** DiodeTransistorPmos: -2.85719e+07 muA
** NormalTransistorPmos: -2.85729e+07 muA
** NormalTransistorPmos: -2.85719e+07 muA
** DiodeTransistorPmos: -2.85729e+07 muA
** NormalTransistorNmos: 1.19681e+08 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 6.00477e+08 muA
** NormalTransistorPmos: -6.00476e+08 muA
** DiodeTransistorNmos: 6.25391e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.11331e+08 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.06001  V
** out: 2.5  V
** outFirstStage: 4.12001  V
** outVoltageBiasXXnXX1: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.28001  V
** innerTransistorStack2Load2: 4.28101  V
** out1: 3.56201  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END