** Name: two_stage_single_output_op_amp_51_11

.MACRO two_stage_single_output_op_amp_51_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=28e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=12e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=89e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=5e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=28e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=12e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=60e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=586e-6
mMainBias11 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=24e-6
mSecondStage1StageBias12 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=598e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=4e-6 W=22e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=5e-6 W=189e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=338e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=338e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=5e-6 W=524e-6
mFoldedCascodeFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=5e-6 W=189e-6
mMainBias21 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=308e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.6001e-12
.EOM two_stage_single_output_op_amp_51_11

** Expected Performance Values: 
** Gain: 167 dB
** Power consumption: 4.02901 mW
** Area: 14993 (mu_m)^2
** Transit frequency: 2.60201 MHz
** Transit frequency with error factor: 2.60227 MHz
** Slew rate: 4.60475 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** VoutMax: 4.25 V
** VoutMin: 0.410001 V
** VcmMax: 5.17001 V
** VcmMin: 0.870001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00451e+07 muA
** NormalTransistorNmos: 2.14841e+07 muA
** NormalTransistorPmos: -7.41139e+07 muA
** NormalTransistorPmos: -5.37089e+07 muA
** NormalTransistorPmos: -8.05619e+07 muA
** NormalTransistorPmos: -5.37119e+07 muA
** NormalTransistorPmos: -8.05669e+07 muA
** NormalTransistorNmos: 5.37101e+07 muA
** NormalTransistorNmos: 5.37111e+07 muA
** DiodeTransistorNmos: 5.37101e+07 muA
** NormalTransistorNmos: 5.37091e+07 muA
** NormalTransistorNmos: 2.68541e+07 muA
** NormalTransistorNmos: 2.68541e+07 muA
** NormalTransistorNmos: 5.28963e+08 muA
** NormalTransistorNmos: 5.28962e+08 muA
** NormalTransistorPmos: -5.28962e+08 muA
** NormalTransistorPmos: -5.28961e+08 muA
** DiodeTransistorNmos: 7.41131e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.00459e+07 muA
** DiodeTransistorPmos: -2.14849e+07 muA


** Expected Voltages: 
** ibias: 0.584001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.20401  V
** out: 2.5  V
** outFirstStage: 4.21501  V
** outVoltageBiasXXnXX1: 1.01201  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.740001  V
** out1: 1.48301  V
** sourceGCC1: 4.53101  V
** sourceGCC2: 4.53101  V
** sourceTransconductance: 1.81201  V
** innerStageBias: 0.379001  V
** innerTransconductance: 4.77901  V


.END