** Name: two_stage_single_output_op_amp_52_11

.MACRO two_stage_single_output_op_amp_52_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=210e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=14e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=210e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=45e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=294e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=11e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=114e-6
mMainBias14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=120e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=157e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=157e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=328e-6
mMainBias19 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=233e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=355e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=120e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.20001e-12
.EOM two_stage_single_output_op_amp_52_11

** Expected Performance Values: 
** Gain: 174 dB
** Power consumption: 6.58401 mW
** Area: 9222 (mu_m)^2
** Transit frequency: 7.19701 MHz
** Transit frequency with error factor: 7.1972 MHz
** Slew rate: 5.91496 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.490001 V
** VcmMax: 5.17001 V
** VcmMin: 0.800001 V


** Expected Currents: 
** NormalTransistorNmos: 1.62454e+08 muA
** NormalTransistorNmos: 7.15001e+06 muA
** NormalTransistorPmos: -1.1867e+08 muA
** NormalTransistorPmos: -4.87359e+07 muA
** NormalTransistorPmos: -8.02769e+07 muA
** NormalTransistorPmos: -4.87359e+07 muA
** NormalTransistorPmos: -8.02769e+07 muA
** DiodeTransistorNmos: 4.87351e+07 muA
** NormalTransistorNmos: 4.87351e+07 muA
** NormalTransistorNmos: 4.87351e+07 muA
** NormalTransistorNmos: 6.30811e+07 muA
** NormalTransistorNmos: 3.15401e+07 muA
** NormalTransistorNmos: 3.15401e+07 muA
** NormalTransistorNmos: 8.58062e+08 muA
** NormalTransistorNmos: 8.58061e+08 muA
** NormalTransistorPmos: -8.58061e+08 muA
** NormalTransistorPmos: -8.58062e+08 muA
** DiodeTransistorNmos: 1.18671e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.62453e+08 muA
** DiodeTransistorPmos: -7.15099e+06 muA


** Expected Voltages: 
** ibias: 0.629001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.09201  V
** out: 2.5  V
** outFirstStage: 4.05201  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.19701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.365001  V
** out1: 0.570001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.92501  V
** innerStageBias: 0.424001  V
** innerTransconductance: 4.61601  V


.END