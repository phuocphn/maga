** Name: two_stage_single_output_op_amp_61_8

.MACRO two_stage_single_output_op_amp_61_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=6e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=338e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=9e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=69e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=344e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=344e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSecondStage1StageBias10 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=413e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=69e-6
mMainBias12 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=46e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=328e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=338e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=59e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=59e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=3e-6 W=350e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=583e-6
mFoldedCascodeFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=161e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.6001e-12
.EOM two_stage_single_output_op_amp_61_8

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 4.50701 mW
** Area: 9172 (mu_m)^2
** Transit frequency: 5.97601 MHz
** Transit frequency with error factor: 5.97531 MHz
** Slew rate: 12.9916 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 4.80001 V
** VoutMin: 0.740001 V
** VcmMax: 3.06001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.04591e+07 muA
** NormalTransistorNmos: 1.06751e+07 muA
** NormalTransistorNmos: 1.4898e+08 muA
** NormalTransistorNmos: 2.24972e+08 muA
** NormalTransistorNmos: 1.4898e+08 muA
** NormalTransistorNmos: 2.24972e+08 muA
** DiodeTransistorPmos: -1.48979e+08 muA
** NormalTransistorPmos: -1.48979e+08 muA
** NormalTransistorPmos: -1.48979e+08 muA
** NormalTransistorPmos: -1.51986e+08 muA
** NormalTransistorPmos: -1.51987e+08 muA
** NormalTransistorPmos: -7.59929e+07 muA
** NormalTransistorPmos: -7.59929e+07 muA
** NormalTransistorNmos: 4.00319e+08 muA
** NormalTransistorNmos: 4.00318e+08 muA
** NormalTransistorPmos: -4.00318e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.04599e+07 muA
** DiodeTransistorPmos: -1.06759e+07 muA


** Expected Voltages: 
** ibias: 1.20501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.23901  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.27501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.51901  V
** innerTransistorStack2Load2: 4.64301  V
** out1: 4.27901  V
** sourceGCC1: 0.522001  V
** sourceGCC2: 0.522001  V
** sourceTransconductance: 3.44201  V
** innerStageBias: 0.614001  V


.END