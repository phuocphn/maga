** Name: two_stage_single_output_op_amp_44_1

.MACRO two_stage_single_output_op_amp_44_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=217e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=240e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=240e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=7e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 outInputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=92e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=203e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=203e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=27e-6
mFoldedCascodeFirstStageLoad9 outFirstStage outInputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=92e-6
mFoldedCascodeFirstStageLoad10 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=240e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=9e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=9e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=62e-6
mSecondStage1StageBias14 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=401e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=4e-6 W=240e-6
mMainBias16 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=105e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_44_1

** Expected Performance Values: 
** Gain: 111 dB
** Power consumption: 5.05901 mW
** Area: 7809 (mu_m)^2
** Transit frequency: 4.18901 MHz
** Transit frequency with error factor: 4.18836 MHz
** Slew rate: 18.2851 V/mu_s
** Phase margin: 65.3172°
** CMRR: 127 dB
** VoutMax: 4.51001 V
** VoutMin: 0.510001 V
** VcmMax: 3.20001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.5237e+08 muA
** NormalTransistorNmos: 8.37301e+07 muA
** NormalTransistorNmos: 1.28881e+08 muA
** NormalTransistorNmos: 8.37291e+07 muA
** NormalTransistorNmos: 1.28881e+08 muA
** NormalTransistorPmos: -8.37309e+07 muA
** NormalTransistorPmos: -8.37299e+07 muA
** DiodeTransistorPmos: -8.37309e+07 muA
** NormalTransistorPmos: -9.02999e+07 muA
** NormalTransistorPmos: -4.51499e+07 muA
** NormalTransistorPmos: -4.51499e+07 muA
** NormalTransistorNmos: 5.81683e+08 muA
** NormalTransistorPmos: -5.81682e+08 muA
** DiodeTransistorNmos: 1.52371e+08 muA
** DiodeTransistorNmos: 1.52372e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 3.94401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.912001  V
** outInputVoltageBiasXXnXX1: 1.11701  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.15601  V
** out1: 3.31201  V
** sourceGCC1: 0.532001  V
** sourceGCC2: 0.532001  V
** sourceTransconductance: 3.81001  V


.END