** Name: two_stage_single_output_op_amp_113_11

.MACRO two_stage_single_output_op_amp_113_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=6e-6
mMainBias2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=117e-6
mTelescopicFirstStageLoad4 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=157e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=90e-6
mSecondStage1StageBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mTelescopicFirstStageLoad7 FirstStageYinnerLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=40e-6
mTelescopicFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=265e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=10e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=473e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=136e-6
mMainBias13 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=286e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=497e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=40e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=80e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=503e-6
mSecondStage1Transconductor18 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=565e-6
mTelescopicFirstStageLoad19 outFirstStage FirstStageYinnerLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=157e-6
mMainBias20 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=152e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.80001e-12
.EOM two_stage_single_output_op_amp_113_11

** Expected Performance Values: 
** Gain: 147 dB
** Power consumption: 5.79601 mW
** Area: 10333 (mu_m)^2
** Transit frequency: 5.14801 MHz
** Transit frequency with error factor: 5.14519 MHz
** Slew rate: 16.8431 V/mu_s
** Phase margin: 60.1606°
** CMRR: 88 dB
** VoutMax: 4.47001 V
** VoutMin: 0.710001 V
** VcmMax: 4.47001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorNmos: 1.33812e+08 muA
** NormalTransistorNmos: 2.82039e+08 muA
** NormalTransistorPmos: -2.21863e+08 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorNmos: 2.59959e+08 muA
** NormalTransistorNmos: 2.5996e+08 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 4.73301e+08 muA
** NormalTransistorNmos: 4.733e+08 muA
** NormalTransistorPmos: -4.733e+08 muA
** NormalTransistorPmos: -4.73301e+08 muA
** DiodeTransistorNmos: 2.21864e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.33811e+08 muA
** DiodeTransistorPmos: -2.82038e+08 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.57501  V
** inputVoltageBiasXXpXX1: 1.93601  V
** out: 2.5  V
** outFirstStage: 4.20601  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXnXX1: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerLoad2: 4.21701  V
** innerStageBias: 0.478001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.606001  V
** innerTransconductance: 2.80501  V


.END