** Name: two_stage_single_output_op_amp_118_9

.MACRO two_stage_single_output_op_amp_118_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=6e-6 W=28e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=5e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=25e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=600e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=4e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=127e-6
mMainBias7 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=10e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=42e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=29e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=10e-6 W=97e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=10e-6 W=97e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias13 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=28e-6
mSecondStage1StageBias14 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=600e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=29e-6
mMainBias16 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=185e-6
mTelescopicFirstStageStageBias18 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=25e-6
mTelescopicFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=127e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=466e-6
mTelescopicFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=202e-6
mMainBias22 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=18e-6
mMainBias23 outVoltageBiasXXnXX3 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=20e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.60001e-12
.EOM two_stage_single_output_op_amp_118_9

** Expected Performance Values: 
** Gain: 154 dB
** Power consumption: 1.75501 mW
** Area: 14970 (mu_m)^2
** Transit frequency: 4.05301 MHz
** Transit frequency with error factor: 4.05252 MHz
** Slew rate: 4.859 V/mu_s
** Phase margin: 60.1606°
** CMRR: 151 dB
** VoutMax: 4.84001 V
** VoutMin: 0.720001 V
** VcmMax: 4.29001 V
** VcmMin: 1.47001 V


** Expected Currents: 
** NormalTransistorNmos: 5.04301e+06 muA
** NormalTransistorNmos: 6.62301e+07 muA
** NormalTransistorPmos: -9.22999e+06 muA
** NormalTransistorPmos: -1.00589e+07 muA
** NormalTransistorNmos: 1.84741e+07 muA
** NormalTransistorNmos: 1.84741e+07 muA
** DiodeTransistorPmos: -1.84749e+07 muA
** NormalTransistorPmos: -1.84749e+07 muA
** NormalTransistorPmos: -1.84749e+07 muA
** NormalTransistorNmos: 4.70071e+07 muA
** DiodeTransistorNmos: 4.70061e+07 muA
** NormalTransistorNmos: 1.84751e+07 muA
** NormalTransistorNmos: 1.84751e+07 muA
** NormalTransistorNmos: 2.13455e+08 muA
** DiodeTransistorNmos: 2.13454e+08 muA
** NormalTransistorPmos: -2.13454e+08 muA
** DiodeTransistorNmos: 9.22901e+06 muA
** NormalTransistorNmos: 9.22801e+06 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 1.00581e+07 muA
** DiodeTransistorPmos: -5.04399e+06 muA
** DiodeTransistorPmos: -6.62309e+07 muA


** Expected Voltages: 
** ibias: 1.12701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.27601  V
** outInputVoltageBiasXXnXX1: 1.32401  V
** outSourceVoltageBiasXXnXX1: 0.662001  V
** outSourceVoltageBiasXXnXX2: 0.564001  V
** outVoltageBiasXXnXX3: 2.65001  V
** outVoltageBiasXXpXX0: 3.90301  V
** outVoltageBiasXXpXX1: 3.71201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 4.45101  V
** out1: 4.21401  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.662001  V
** inner: 0.563001  V


.END