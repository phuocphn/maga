** Name: two_stage_single_output_op_amp_134_5

.MACRO two_stage_single_output_op_amp_134_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=9e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=27e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=4e-6 W=27e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=18e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=8e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=349e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=191e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=191e-6
mSimpleFirstStageLoad10 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=58e-6
mMainBias11 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=25e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=363e-6
mSimpleFirstStageLoad13 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=58e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=22e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=27e-6
mSimpleFirstStageTransconductor16 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=45e-6
mSimpleFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=126e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=8e-6
mSecondStage1StageBias19 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=349e-6
mSimpleFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=27e-6
mSimpleFirstStageTransconductor21 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=45e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_134_5

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 4.54901 mW
** Area: 10266 (mu_m)^2
** Transit frequency: 5.20101 MHz
** Transit frequency with error factor: 5.18644 MHz
** Slew rate: 24.6309 V/mu_s
** Phase margin: 60.1606°
** CMRR: 80 dB
** VoutMax: 3.02001 V
** VoutMin: 0.380001 V
** VcmMax: 3.01001 V
** VcmMin: -0.129999 V


** Expected Currents: 
** NormalTransistorNmos: 1.43881e+07 muA
** NormalTransistorNmos: 1.63501e+07 muA
** DiodeTransistorPmos: -6.85349e+07 muA
** DiodeTransistorPmos: -6.85349e+07 muA
** NormalTransistorPmos: -6.85349e+07 muA
** NormalTransistorPmos: -6.85349e+07 muA
** NormalTransistorNmos: 1.25647e+08 muA
** NormalTransistorNmos: 1.25646e+08 muA
** NormalTransistorNmos: 1.25647e+08 muA
** NormalTransistorNmos: 1.25646e+08 muA
** NormalTransistorPmos: -1.14224e+08 muA
** NormalTransistorPmos: -5.71119e+07 muA
** NormalTransistorPmos: -5.71119e+07 muA
** NormalTransistorNmos: 6.17729e+08 muA
** NormalTransistorPmos: -6.17728e+08 muA
** DiodeTransistorPmos: -6.17729e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.43889e+07 muA
** NormalTransistorPmos: -1.43899e+07 muA
** DiodeTransistorPmos: -1.63509e+07 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.75701  V
** out: 2.5  V
** outFirstStage: 0.782001  V
** outInputVoltageBiasXXpXX1: 2.45801  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 3.72901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.478001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.478001  V
** out1: 2.37201  V
** sourceTransconductance: 3.81401  V
** inner: 3.72801  V


.END