** Name: two_stage_single_output_op_amp_19_6

.MACRO two_stage_single_output_op_amp_19_6 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=97e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=53e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=25e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=250e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=97e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=599e-6
mSecondStage1Transconductor10 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=50e-6
mMainBias12 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=288e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=178e-6
mSimpleFirstStageStageBias14 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=387e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mSecondStage1StageBias17 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=250e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=178e-6
mMainBias19 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=35e-6
mMainBias20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=182e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.8001e-12
.EOM two_stage_single_output_op_amp_19_6

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 14.7191 mW
** Area: 5629 (mu_m)^2
** Transit frequency: 28.8491 MHz
** Transit frequency with error factor: 28.8118 MHz
** Slew rate: 56.0518 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** negPSRR: 100 dB
** posPSRR: 142 dB
** VoutMax: 3.12001 V
** VoutMin: 0.390001 V
** VcmMax: 3.03001 V
** VcmMin: 0.300001 V


** Expected Currents: 
** NormalTransistorNmos: 1.94194e+08 muA
** NormalTransistorPmos: -3.54849e+07 muA
** NormalTransistorPmos: -1.80928e+08 muA
** DiodeTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorPmos: -6.08327e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorNmos: 1.90491e+09 muA
** NormalTransistorNmos: 1.90491e+09 muA
** NormalTransistorPmos: -1.9049e+09 muA
** DiodeTransistorPmos: -1.90491e+09 muA
** DiodeTransistorNmos: 3.54841e+07 muA
** DiodeTransistorNmos: 1.80929e+08 muA
** DiodeTransistorPmos: -1.94193e+08 muA
** NormalTransistorPmos: -1.94193e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.598001  V
** outInputVoltageBiasXXpXX1: 2.56001  V
** outSourceVoltageBiasXXpXX1: 3.78001  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.623001  V
** outVoltageBiasXXnXX1: 0.865001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.598001  V
** innerStageBias: 4.25801  V
** innerTransistorStack2Load1: 0.193001  V
** sourceTransconductance: 3.37201  V
** innerTransconductance: 0.266001  V
** inner: 3.78001  V


.END