** Name: two_stage_single_output_op_amp_64_8

.MACRO two_stage_single_output_op_amp_64_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=20e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=21e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=47e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=8e-6 W=152e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=384e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 outInputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=314e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=158e-6
mFoldedCascodeFirstStageLoad12 outFirstStage outInputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=29e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=8e-6 W=384e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=152e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=118e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=47e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=600e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_64_8

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 3.67601 mW
** Area: 14531 (mu_m)^2
** Transit frequency: 3.30401 MHz
** Transit frequency with error factor: 3.30411 MHz
** Slew rate: 5.6194 V/mu_s
** Phase margin: 64.1713°
** CMRR: 141 dB
** VoutMax: 4.25 V
** VoutMin: 0.770001 V
** VcmMax: 3.26001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -3.99979e+07 muA
** NormalTransistorNmos: 2.53751e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorNmos: 2.53751e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** DiodeTransistorPmos: -2.53759e+07 muA
** DiodeTransistorPmos: -2.53769e+07 muA
** NormalTransistorPmos: -2.53759e+07 muA
** NormalTransistorPmos: -2.53769e+07 muA
** NormalTransistorPmos: -2.54389e+07 muA
** DiodeTransistorPmos: -2.54399e+07 muA
** NormalTransistorPmos: -1.27189e+07 muA
** NormalTransistorPmos: -1.27189e+07 muA
** NormalTransistorNmos: 5.99051e+08 muA
** NormalTransistorNmos: 5.9905e+08 muA
** NormalTransistorPmos: -5.9905e+08 muA
** DiodeTransistorNmos: 3.99971e+07 muA
** DiodeTransistorNmos: 3.99981e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.52701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.11301  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.26401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.24501  V
** innerTransistorStack2Load2: 4.24401  V
** out1: 3.50701  V
** sourceGCC1: 0.534001  V
** sourceGCC2: 0.534001  V
** sourceTransconductance: 3.33401  V
** innerStageBias: 0.496001  V
** inner: 4.26201  V


.END