** Name: two_stage_single_output_op_amp_4_5

.MACRO two_stage_single_output_op_amp_4_5 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=30e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=30e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=16e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=9e-6 W=195e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=7e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=447e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=30e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=357e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=30e-6
mMainBias10 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=45e-6
mSimpleFirstStageTransconductor11 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=71e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=9e-6 W=446e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=7e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=447e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=71e-6
mMainBias16 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=9e-6 W=75e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_4_5

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 3.75501 mW
** Area: 14834 (mu_m)^2
** Transit frequency: 4.92301 MHz
** Transit frequency with error factor: 4.92069 MHz
** Slew rate: 5.12091 V/mu_s
** Phase margin: 76.2034°
** CMRR: 106 dB
** negPSRR: 101 dB
** posPSRR: 106 dB
** VoutMax: 3 V
** VoutMin: 0.300001 V
** VcmMax: 4.11001 V
** VcmMin: 0.550001 V


** Expected Currents: 
** NormalTransistorNmos: 1.07501e+07 muA
** NormalTransistorPmos: -3.89899e+06 muA
** DiodeTransistorNmos: 1.15921e+07 muA
** DiodeTransistorNmos: 1.15911e+07 muA
** NormalTransistorNmos: 1.15921e+07 muA
** NormalTransistorNmos: 1.15911e+07 muA
** NormalTransistorPmos: -2.31859e+07 muA
** NormalTransistorPmos: -1.15929e+07 muA
** NormalTransistorPmos: -1.15929e+07 muA
** NormalTransistorNmos: 6.93257e+08 muA
** NormalTransistorPmos: -6.93256e+08 muA
** DiodeTransistorPmos: -6.93256e+08 muA
** DiodeTransistorNmos: 3.89801e+06 muA
** DiodeTransistorPmos: -1.07509e+07 muA
** NormalTransistorPmos: -1.07519e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.707001  V
** outInputVoltageBiasXXpXX1: 2.43601  V
** outSourceVoltageBiasXXpXX1: 3.71801  V
** outVoltageBiasXXnXX0: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 1.11201  V
** innerSourceLoad1: 0.556001  V
** innerTransistorStack2Load1: 0.556001  V
** sourceTransconductance: 3.22901  V
** inner: 3.71501  V


.END