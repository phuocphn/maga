** Name: two_stage_single_output_op_amp_32_11

.MACRO two_stage_single_output_op_amp_32_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=10e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=264e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=218e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=50e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=12e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=528e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=264e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=301e-6
mSecondStage1StageBias13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=552e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=50e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=445e-6
mSimpleFirstStageLoad16 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=508e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=424e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=48e-6
mMainBias20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=437e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.80001e-12
.EOM two_stage_single_output_op_amp_32_11

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 9.43001 mW
** Area: 10996 (mu_m)^2
** Transit frequency: 4.95401 MHz
** Transit frequency with error factor: 4.95098 MHz
** Slew rate: 4.66924 V/mu_s
** Phase margin: 60.1606°
** CMRR: 104 dB
** negPSRR: 117 dB
** posPSRR: 103 dB
** VoutMax: 4.25 V
** VoutMin: 0.710001 V
** VcmMax: 4.36001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 2.98632e+08 muA
** NormalTransistorNmos: 4.36596e+08 muA
** NormalTransistorPmos: -5.87875e+08 muA
** NormalTransistorPmos: -1.36059e+07 muA
** NormalTransistorPmos: -1.36059e+07 muA
** DiodeTransistorPmos: -1.36059e+07 muA
** NormalTransistorNmos: 2.72091e+07 muA
** DiodeTransistorNmos: 2.72081e+07 muA
** NormalTransistorNmos: 1.36051e+07 muA
** NormalTransistorNmos: 1.36051e+07 muA
** NormalTransistorNmos: 5.25678e+08 muA
** NormalTransistorNmos: 5.25677e+08 muA
** NormalTransistorPmos: -5.25677e+08 muA
** NormalTransistorPmos: -5.25678e+08 muA
** DiodeTransistorNmos: 5.87876e+08 muA
** NormalTransistorNmos: 5.87876e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.98631e+08 muA
** DiodeTransistorPmos: -4.36595e+08 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.82001  V
** out: 2.5  V
** outFirstStage: 3.95301  V
** outInputVoltageBiasXXnXX1: 1.13601  V
** outSourceVoltageBiasXXnXX1: 0.568001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.23501  V
** out1: 3.38901  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.561001  V
** innerTransconductance: 4.51301  V
** inner: 0.568001  V


.END