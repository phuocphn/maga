** Name: two_stage_single_output_op_amp_71_11

.MACRO two_stage_single_output_op_amp_71_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=19e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=10e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=108e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=312e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=26e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=26e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=9e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=564e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=553e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=588e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=19e-6
mMainBias14 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=36e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerLoad2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=76e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=211e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=211e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=556e-6
mSecondStage1Transconductor19 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=496e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=76e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_71_11

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 6.01001 mW
** Area: 12184 (mu_m)^2
** Transit frequency: 3.17501 MHz
** Transit frequency with error factor: 3.17273 MHz
** Slew rate: 3.5002 V/mu_s
** Phase margin: 71.6198°
** CMRR: 102 dB
** VoutMax: 4.31001 V
** VoutMin: 0.710001 V
** VcmMax: 5.19001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 5.48284e+08 muA
** NormalTransistorNmos: 3.54051e+07 muA
** NormalTransistorPmos: -1.58469e+07 muA
** NormalTransistorPmos: -2.41859e+07 muA
** NormalTransistorPmos: -1.58469e+07 muA
** NormalTransistorPmos: -2.41859e+07 muA
** DiodeTransistorNmos: 1.58461e+07 muA
** NormalTransistorNmos: 1.58461e+07 muA
** NormalTransistorNmos: 1.66761e+07 muA
** NormalTransistorNmos: 1.66771e+07 muA
** NormalTransistorNmos: 8.33801e+06 muA
** NormalTransistorNmos: 8.33801e+06 muA
** NormalTransistorNmos: 5.59961e+08 muA
** NormalTransistorNmos: 5.5996e+08 muA
** NormalTransistorPmos: -5.5996e+08 muA
** NormalTransistorPmos: -5.59961e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.48283e+08 muA
** DiodeTransistorPmos: -3.54059e+07 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.09901  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX2: 4.22501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.718001  V
** innerStageBias: 0.501001  V
** sourceGCC1: 4.40201  V
** sourceGCC2: 4.40201  V
** sourceTransconductance: 1.91001  V
** innerStageBias: 0.561001  V
** innerTransconductance: 4.60401  V


.END