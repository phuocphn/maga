** Name: two_stage_single_output_op_amp_61_11

.MACRO two_stage_single_output_op_amp_61_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=15e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=7e-6 W=269e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=13e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=23e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=45e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=45e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=170e-6
mSecondStage1StageBias11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=301e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=23e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=101e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=7e-6 W=269e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=86e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=86e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=23e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=448e-6
mSecondStage1Transconductor20 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=140e-6
mFoldedCascodeFirstStageLoad21 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=41e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_61_11

** Expected Performance Values: 
** Gain: 177 dB
** Power consumption: 2.91701 mW
** Area: 10314 (mu_m)^2
** Transit frequency: 4.36201 MHz
** Transit frequency with error factor: 4.36237 MHz
** Slew rate: 4.30673 V/mu_s
** Phase margin: 64.7443°
** CMRR: 146 dB
** VoutMax: 4.28001 V
** VoutMin: 0.780001 V
** VcmMax: 3.17001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.11687e+08 muA
** NormalTransistorNmos: 2.61901e+06 muA
** NormalTransistorNmos: 1.94551e+07 muA
** NormalTransistorNmos: 2.94301e+07 muA
** NormalTransistorNmos: 1.94551e+07 muA
** NormalTransistorNmos: 2.94301e+07 muA
** DiodeTransistorPmos: -1.94559e+07 muA
** NormalTransistorPmos: -1.94559e+07 muA
** NormalTransistorPmos: -1.94559e+07 muA
** NormalTransistorPmos: -1.99529e+07 muA
** NormalTransistorPmos: -1.99539e+07 muA
** NormalTransistorPmos: -9.97599e+06 muA
** NormalTransistorPmos: -9.97599e+06 muA
** NormalTransistorNmos: 4.00319e+08 muA
** NormalTransistorNmos: 4.00318e+08 muA
** NormalTransistorPmos: -4.00318e+08 muA
** NormalTransistorPmos: -4.00319e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.11686e+08 muA
** DiodeTransistorPmos: -2.61999e+06 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.11901  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX2: 4.11901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.47001  V
** innerTransistorStack2Load2: 4.41301  V
** out1: 4.26701  V
** sourceGCC1: 0.537001  V
** sourceGCC2: 0.537001  V
** sourceTransconductance: 3.22501  V
** innerStageBias: 0.493001  V
** innerTransconductance: 4.64901  V


.END