** Name: two_stage_single_output_op_amp_11_12

.MACRO two_stage_single_output_op_amp_11_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=5e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=142e-6
mSimpleFirstStageLoad4 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=437e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=223e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=11e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=280e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=145e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=142e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=280e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=17e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=159e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=223e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=556e-6
mSecondStage1Transconductor17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad18 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=437e-6
mMainBias19 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=41e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.1001e-12
.EOM two_stage_single_output_op_amp_11_12

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 8.92301 mW
** Area: 12708 (mu_m)^2
** Transit frequency: 11.1161 MHz
** Transit frequency with error factor: 11.1105 MHz
** Slew rate: 10.4768 V/mu_s
** Phase margin: 60.1606°
** CMRR: 110 dB
** negPSRR: 107 dB
** posPSRR: 100 dB
** VoutMax: 4.25 V
** VoutMin: 1.79001 V
** VcmMax: 3.92001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorNmos: 1.39721e+07 muA
** NormalTransistorNmos: 1.31994e+08 muA
** NormalTransistorPmos: -5.14789e+07 muA
** DiodeTransistorPmos: -5.92569e+07 muA
** DiodeTransistorPmos: -5.92579e+07 muA
** NormalTransistorPmos: -5.92569e+07 muA
** NormalTransistorPmos: -5.92579e+07 muA
** NormalTransistorNmos: 1.18512e+08 muA
** NormalTransistorNmos: 5.92561e+07 muA
** NormalTransistorNmos: 5.92561e+07 muA
** NormalTransistorNmos: 1.45873e+09 muA
** DiodeTransistorNmos: 1.45873e+09 muA
** NormalTransistorPmos: -1.45872e+09 muA
** NormalTransistorPmos: -1.45872e+09 muA
** DiodeTransistorNmos: 5.14781e+07 muA
** NormalTransistorNmos: 5.14771e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.39729e+07 muA
** DiodeTransistorPmos: -1.31993e+08 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.05301  V
** outInputVoltageBiasXXnXX1: 2.19801  V
** outSourceVoltageBiasXXnXX1: 1.09901  V
** outVoltageBiasXXpXX0: 3.73201  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.51001  V
** innerSourceLoad1: 4.22501  V
** innerTransistorStack2Load1: 4.22501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.61701  V
** inner: 1.09301  V


.END