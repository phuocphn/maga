** Name: two_stage_single_output_op_amp_54_12

.MACRO two_stage_single_output_op_amp_54_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=14e-6
mMainBias2 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=8e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=384e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=26e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=308e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=72e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=72e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=40e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=384e-6
mFoldedCascodeFirstStageLoad15 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=308e-6
mMainBias16 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=14e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=438e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=353e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=353e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=461e-6
mMainBias21 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=151e-6
mMainBias22 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=63e-6
mSecondStage1Transconductor23 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad24 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=438e-6
mMainBias25 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.6001e-12
.EOM two_stage_single_output_op_amp_54_12

** Expected Performance Values: 
** Gain: 172 dB
** Power consumption: 6.80601 mW
** Area: 14969 (mu_m)^2
** Transit frequency: 4.79401 MHz
** Transit frequency with error factor: 4.79407 MHz
** Slew rate: 6.01104 V/mu_s
** Phase margin: 60.1606°
** CMRR: 139 dB
** VoutMax: 4.25 V
** VoutMin: 0.990001 V
** VcmMax: 5.20001 V
** VcmMin: 1.16001 V


** Expected Currents: 
** NormalTransistorNmos: 3.49061e+07 muA
** NormalTransistorPmos: -1.94429e+07 muA
** NormalTransistorPmos: -5.85259e+07 muA
** NormalTransistorPmos: -2.44409e+07 muA
** NormalTransistorPmos: -8.89429e+07 muA
** NormalTransistorPmos: -1.37834e+08 muA
** NormalTransistorPmos: -8.89429e+07 muA
** NormalTransistorPmos: -1.37834e+08 muA
** NormalTransistorNmos: 8.89421e+07 muA
** NormalTransistorNmos: 8.89411e+07 muA
** NormalTransistorNmos: 8.89421e+07 muA
** NormalTransistorNmos: 8.89411e+07 muA
** NormalTransistorNmos: 9.77811e+07 muA
** NormalTransistorNmos: 4.88911e+07 muA
** NormalTransistorNmos: 4.88911e+07 muA
** NormalTransistorNmos: 9.28135e+08 muA
** DiodeTransistorNmos: 9.28134e+08 muA
** NormalTransistorPmos: -9.28134e+08 muA
** NormalTransistorPmos: -9.28135e+08 muA
** DiodeTransistorNmos: 1.94421e+07 muA
** NormalTransistorNmos: 1.94411e+07 muA
** DiodeTransistorNmos: 5.85251e+07 muA
** DiodeTransistorNmos: 2.44401e+07 muA
** DiodeTransistorPmos: -3.49069e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.22801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.07501  V
** inputVoltageBiasXXnXX3: 0.945001  V
** out: 2.5  V
** outFirstStage: 4.10001  V
** outInputVoltageBiasXXnXX1: 1.39401  V
** outSourceVoltageBiasXXnXX1: 0.697001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.700001  V
** innerTransistorStack1Load2: 0.494001  V
** innerTransistorStack2Load2: 0.495001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.875  V
** innerTransconductance: 4.66401  V
** inner: 0.695001  V


.END