** Name: two_stage_single_output_op_amp_118_10

.MACRO two_stage_single_output_op_amp_118_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=13e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=12e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=49e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=10e-6 W=12e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=104e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=9e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=10e-6 W=61e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=49e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=49e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=12e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=10e-6 W=61e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=165e-6
mTelescopicFirstStageStageBias16 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=49e-6
mTelescopicFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=104e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=347e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mTelescopicFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=29e-6
mMainBias21 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=13e-6
mMainBias22 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=15e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_118_10

** Expected Performance Values: 
** Gain: 152 dB
** Power consumption: 3.23501 mW
** Area: 9383 (mu_m)^2
** Transit frequency: 2.68401 MHz
** Transit frequency with error factor: 2.6838 MHz
** Slew rate: 3.51066 V/mu_s
** Phase margin: 60.1606°
** CMRR: 154 dB
** VoutMax: 4.52001 V
** VoutMin: 0.210001 V
** VcmMax: 4.38001 V
** VcmMin: 1.52001 V


** Expected Currents: 
** NormalTransistorNmos: 5.43001e+06 muA
** NormalTransistorNmos: 1.27061e+08 muA
** NormalTransistorPmos: -7.82999e+06 muA
** NormalTransistorPmos: -9.05299e+06 muA
** NormalTransistorNmos: 1.16661e+07 muA
** NormalTransistorNmos: 1.16651e+07 muA
** DiodeTransistorPmos: -1.16669e+07 muA
** NormalTransistorPmos: -1.16659e+07 muA
** NormalTransistorPmos: -1.16669e+07 muA
** NormalTransistorNmos: 3.23831e+07 muA
** DiodeTransistorNmos: 3.23821e+07 muA
** NormalTransistorNmos: 1.16661e+07 muA
** NormalTransistorNmos: 1.16661e+07 muA
** NormalTransistorNmos: 4.64299e+08 muA
** NormalTransistorPmos: -4.64298e+08 muA
** NormalTransistorPmos: -4.64299e+08 muA
** DiodeTransistorNmos: 7.82901e+06 muA
** NormalTransistorNmos: 7.82901e+06 muA
** DiodeTransistorNmos: 9.05201e+06 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.43099e+06 muA
** DiodeTransistorPmos: -1.2706e+08 muA


** Expected Voltages: 
** ibias: 0.618001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.16101  V
** outInputVoltageBiasXXnXX1: 1.36801  V
** outSourceVoltageBiasXXnXX1: 0.684001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 3.91501  V
** outVoltageBiasXXpXX1: 3.59701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 4.31101  V
** out1: 4.27701  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.36901  V
** inner: 0.684001  V


.END