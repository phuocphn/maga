** Name: two_stage_single_output_op_amp_206_8

.MACRO two_stage_single_output_op_amp_206_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=8e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=6e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=89e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=37e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=114e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=13e-6
mSimpleFirstStageTransconductor9 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=13e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=37e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=107e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=89e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=6e-6 W=103e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=8e-6 W=10e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=13e-6
mSimpleFirstStageLoad17 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=7e-6 W=264e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=60e-6
mSimpleFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=60e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=58e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=574e-6
mSimpleFirstStageLoad22 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=264e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_206_8

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 5.11601 mW
** Area: 14011 (mu_m)^2
** Transit frequency: 3.26001 MHz
** Transit frequency with error factor: 3.25841 MHz
** Slew rate: 3.50015 V/mu_s
** Phase margin: 64.7443°
** CMRR: 110 dB
** VoutMax: 4.25 V
** VoutMin: 1.89001 V
** VcmMax: 4.59001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorPmos: -3.88159e+07 muA
** NormalTransistorPmos: -4.54009e+07 muA
** DiodeTransistorNmos: 3.85991e+07 muA
** NormalTransistorNmos: 3.86001e+07 muA
** NormalTransistorNmos: 3.86011e+07 muA
** DiodeTransistorNmos: 3.86001e+07 muA
** NormalTransistorPmos: -4.66329e+07 muA
** NormalTransistorPmos: -4.66339e+07 muA
** NormalTransistorPmos: -4.66349e+07 muA
** NormalTransistorPmos: -4.66339e+07 muA
** NormalTransistorNmos: 1.60661e+07 muA
** DiodeTransistorNmos: 1.60651e+07 muA
** NormalTransistorNmos: 8.03301e+06 muA
** NormalTransistorNmos: 8.03301e+06 muA
** NormalTransistorNmos: 8.25659e+08 muA
** NormalTransistorNmos: 8.25658e+08 muA
** NormalTransistorPmos: -8.25658e+08 muA
** DiodeTransistorNmos: 3.88151e+07 muA
** NormalTransistorNmos: 3.88141e+07 muA
** DiodeTransistorNmos: 4.54001e+07 muA
** DiodeTransistorNmos: 4.54011e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 2.27501  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.21401  V
** outSourceVoltageBiasXXnXX1: 0.607001  V
** outSourceVoltageBiasXXnXX2: 1.14101  V
** outSourceVoltageBiasXXpXX1: 3.88501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.08301  V
** innerTransistorStack1Load1: 1.08401  V
** innerTransistorStack1Load2: 3.96101  V
** innerTransistorStack2Load2: 3.96101  V
** sourceTransconductance: 1.92401  V
** innerStageBias: 1.12001  V
** inner: 0.605001  V


.END