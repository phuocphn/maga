** Name: symmetrical_op_amp142

.MACRO symmetrical_op_amp142 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=11e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=11e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=117e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=114e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=10e-6 W=12e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=54e-6
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=54e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=121e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=121e-6
mSymmetricalFirstStageLoad10 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=85e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=7e-6 W=86e-6
mSecondStage1Transconductor12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=7e-6 W=86e-6
mSymmetricalFirstStageLoad13 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=85e-6
mMainBias14 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=27e-6
mSymmetricalFirstStageStageBias15 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=600e-6
mSymmetricalFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=10e-6 W=108e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=114e-6
mSymmetricalFirstStageTransconductor18 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=55e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=10e-6 W=104e-6
mSymmetricalFirstStageTransconductor20 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=55e-6
mMainBias21 out2FirstStage ibias sourcePmos sourcePmos pmos4 L=7e-6 W=227e-6
mMainBias22 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=56e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp142

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 1.11701 mW
** Area: 13715 (mu_m)^2
** Transit frequency: 5.67901 MHz
** Transit frequency with error factor: 5.67934 MHz
** Slew rate: 5.75003 V/mu_s
** Phase margin: 61.3065°
** CMRR: 145 dB
** negPSRR: 50 dB
** posPSRR: 58 dB
** VoutMax: 4.28001 V
** VoutMin: 0.380001 V
** VcmMax: 3.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.20311e+07 muA
** NormalTransistorPmos: -4.83499e+06 muA
** NormalTransistorPmos: -1.95229e+07 muA
** NormalTransistorNmos: 2.59061e+07 muA
** NormalTransistorNmos: 2.59051e+07 muA
** NormalTransistorNmos: 2.59061e+07 muA
** NormalTransistorNmos: 2.59051e+07 muA
** NormalTransistorPmos: -5.18139e+07 muA
** NormalTransistorPmos: -5.18129e+07 muA
** NormalTransistorPmos: -2.59069e+07 muA
** NormalTransistorPmos: -2.59069e+07 muA
** NormalTransistorNmos: 5.76141e+07 muA
** NormalTransistorNmos: 5.76151e+07 muA
** NormalTransistorPmos: -5.76149e+07 muA
** NormalTransistorPmos: -5.76159e+07 muA
** DiodeTransistorPmos: -5.76149e+07 muA
** NormalTransistorNmos: 5.76141e+07 muA
** NormalTransistorNmos: 5.76151e+07 muA
** DiodeTransistorNmos: 4.83401e+06 muA
** DiodeTransistorNmos: 1.95221e+07 muA
** DiodeTransistorPmos: -1.20319e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25301  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 4.26701  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.790001  V
** outVoltageBiasXXnXX0: 0.596001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.76601  V
** innerTransistorStack1Load1: 0.226001  V
** innerTransistorStack2Load1: 0.226001  V
** sourceTransconductance: 3.22601  V
** innerStageBias: 4.80401  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END