** Name: two_stage_single_output_op_amp_148_7

.MACRO two_stage_single_output_op_amp_148_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=23e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=10e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=268e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=154e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=11e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=46e-6
mMainBias9 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=120e-6
mSecondStage1StageBias10 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=23e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=11e-6
mSimpleFirstStageLoad13 FirstStageYinnerOutputLoad1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=261e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=275e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=275e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=392e-6
mSimpleFirstStageLoad17 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=261e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.4001e-12
.EOM two_stage_single_output_op_amp_148_7

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 5.74301 mW
** Area: 6390 (mu_m)^2
** Transit frequency: 4.39901 MHz
** Transit frequency with error factor: 4.39652 MHz
** Slew rate: 4.30416 V/mu_s
** Phase margin: 60.1606°
** CMRR: 116 dB
** VoutMax: 4.58001 V
** VoutMin: 0.240001 V
** VcmMax: 4.99001 V
** VcmMin: 0.800001 V


** Expected Currents: 
** NormalTransistorNmos: 1.19111e+08 muA
** DiodeTransistorNmos: 1.86678e+08 muA
** DiodeTransistorNmos: 1.86677e+08 muA
** NormalTransistorNmos: 1.86676e+08 muA
** NormalTransistorNmos: 1.86677e+08 muA
** NormalTransistorPmos: -2.09255e+08 muA
** NormalTransistorPmos: -2.09254e+08 muA
** NormalTransistorPmos: -2.09253e+08 muA
** NormalTransistorPmos: -2.09254e+08 muA
** NormalTransistorNmos: 4.51571e+07 muA
** NormalTransistorNmos: 2.25781e+07 muA
** NormalTransistorNmos: 2.25781e+07 muA
** NormalTransistorNmos: 6.00903e+08 muA
** NormalTransistorPmos: -6.00902e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.1911e+08 muA
** DiodeTransistorPmos: -1.19109e+08 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.50701  V
** out: 2.5  V
** outFirstStage: 4.02001  V
** outSourceVoltageBiasXXpXX1: 4.22901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerTransistorStack1Load1: 1.15101  V
** innerTransistorStack1Load2: 4.28201  V
** innerTransistorStack2Load1: 1.15201  V
** innerTransistorStack2Load2: 4.28201  V
** sourceTransconductance: 1.93901  V


.END