** Name: two_stage_single_output_op_amp_144_11

.MACRO two_stage_single_output_op_amp_144_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=122e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=25e-6
mSimpleFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=122e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=56e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=331e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=120e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=25e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=28e-6
mMainBias14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=72e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
mSimpleFirstStageLoad17 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=564e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=325e-6
mMainBias19 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=544e-6
mSimpleFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=564e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.9001e-12
.EOM two_stage_single_output_op_amp_144_11

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 14.7471 mW
** Area: 11326 (mu_m)^2
** Transit frequency: 5.47201 MHz
** Transit frequency with error factor: 5.46807 MHz
** Slew rate: 6.19588 V/mu_s
** Phase margin: 60.1606°
** CMRR: 123 dB
** VoutMax: 4.25 V
** VoutMin: 0.570001 V
** VcmMax: 4.66001 V
** VcmMin: 0.830001 V


** Expected Currents: 
** NormalTransistorNmos: 3.50521e+07 muA
** NormalTransistorNmos: 8.95781e+07 muA
** NormalTransistorPmos: -7.63969e+07 muA
** NormalTransistorNmos: 9.59565e+08 muA
** NormalTransistorNmos: 9.59564e+08 muA
** DiodeTransistorNmos: 9.59565e+08 muA
** NormalTransistorPmos: -9.93923e+08 muA
** NormalTransistorPmos: -9.93923e+08 muA
** NormalTransistorPmos: -9.93922e+08 muA
** NormalTransistorPmos: -9.93923e+08 muA
** NormalTransistorNmos: 6.87181e+07 muA
** NormalTransistorNmos: 3.43591e+07 muA
** NormalTransistorNmos: 3.43591e+07 muA
** NormalTransistorNmos: 7.50605e+08 muA
** NormalTransistorNmos: 7.50604e+08 muA
** NormalTransistorPmos: -7.50604e+08 muA
** NormalTransistorPmos: -7.50605e+08 muA
** DiodeTransistorNmos: 7.63961e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.50529e+07 muA
** DiodeTransistorPmos: -8.95789e+07 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.975001  V
** out: 2.5  V
** outFirstStage: 4.07701  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.13001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack1Load2: 4.69201  V
** innerTransistorStack2Load2: 4.69201  V
** out1: 2.09501  V
** sourceTransconductance: 1.91401  V
** innerStageBias: 0.242001  V
** innerTransconductance: 4.64101  V


.END