** Name: two_stage_single_output_op_amp_162_6

.MACRO two_stage_single_output_op_amp_162_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mMainBias4 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=4e-6 W=21e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=211e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=103e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=509e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=170e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=170e-6
mSimpleFirstStageLoad10 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=85e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=129e-6
mSecondStage1Transconductor12 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=389e-6
mSimpleFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=85e-6
mMainBias14 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=390e-6
mSimpleFirstStageTransconductor15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=304e-6
mSimpleFirstStageLoad16 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mSimpleFirstStageStageBias17 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=103e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=211e-6
mMainBias19 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=21e-6
mMainBias20 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=21e-6
mMainBias21 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSecondStage1StageBias22 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=4e-6 W=509e-6
mSimpleFirstStageLoad23 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=12e-6
mSimpleFirstStageTransconductor24 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=304e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.3001e-12
.EOM two_stage_single_output_op_amp_162_6

** Expected Performance Values: 
** Gain: 149 dB
** Power consumption: 2.55501 mW
** Area: 14970 (mu_m)^2
** Transit frequency: 3.64201 MHz
** Transit frequency with error factor: 3.63995 MHz
** Slew rate: 4.16281 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 3.78001 V
** VoutMin: 0.300001 V
** VcmMax: 3.33001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 1.23802e+08 muA
** NormalTransistorPmos: -1.01949e+07 muA
** NormalTransistorPmos: -1.90599e+06 muA
** NormalTransistorPmos: -2.40099e+07 muA
** NormalTransistorPmos: -2.40089e+07 muA
** DiodeTransistorPmos: -2.40099e+07 muA
** NormalTransistorNmos: 5.39661e+07 muA
** NormalTransistorNmos: 5.39651e+07 muA
** NormalTransistorNmos: 5.39651e+07 muA
** NormalTransistorNmos: 5.39651e+07 muA
** NormalTransistorPmos: -5.99149e+07 muA
** DiodeTransistorPmos: -5.99159e+07 muA
** NormalTransistorPmos: -2.99569e+07 muA
** NormalTransistorPmos: -2.99569e+07 muA
** NormalTransistorNmos: 2.47113e+08 muA
** NormalTransistorNmos: 2.47112e+08 muA
** NormalTransistorPmos: -2.47112e+08 muA
** DiodeTransistorPmos: -2.47111e+08 muA
** DiodeTransistorNmos: 1.01941e+07 muA
** DiodeTransistorNmos: 1.90501e+06 muA
** DiodeTransistorPmos: -1.23801e+08 muA
** NormalTransistorPmos: -1.23802e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.21301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.51001  V
** outSourceVoltageBiasXXpXX1: 4.25501  V
** outSourceVoltageBiasXXpXX2: 4.10801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.22401  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 2.91001  V
** sourceTransconductance: 3.24501  V
** innerTransconductance: 0.150001  V
** inner: 4.25501  V
** inner: 4.10201  V


.END