** Name: two_stage_single_output_op_amp_80_11

.MACRO two_stage_single_output_op_amp_80_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
mMainBias2 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=71e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=23e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=223e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=38e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=123e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=33e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=33e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=30e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=30e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=223e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=599e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=23e-6
mSecondStage1StageBias15 out inputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=547e-6
mFoldedCascodeFirstStageLoad16 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=123e-6
mMainBias17 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=44e-6
mFoldedCascodeFirstStageLoad18 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=61e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=525e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=525e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=485e-6
mMainBias22 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=594e-6
mMainBias23 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=596e-6
mSecondStage1Transconductor24 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad25 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=61e-6
mMainBias26 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=45e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.2001e-12
.EOM two_stage_single_output_op_amp_80_11

** Expected Performance Values: 
** Gain: 171 dB
** Power consumption: 10.4171 mW
** Area: 14987 (mu_m)^2
** Transit frequency: 7.46601 MHz
** Transit frequency with error factor: 7.46561 MHz
** Slew rate: 5.11264 V/mu_s
** Phase margin: 60.1606°
** CMRR: 137 dB
** VoutMax: 4.25 V
** VoutMin: 0.5 V
** VcmMax: 5.23001 V
** VcmMin: 1.45001 V


** Expected Currents: 
** NormalTransistorNmos: 9.99581e+07 muA
** NormalTransistorPmos: -1.2e+07 muA
** NormalTransistorPmos: -1.5577e+08 muA
** NormalTransistorPmos: -1.58103e+08 muA
** NormalTransistorPmos: -8.30359e+07 muA
** NormalTransistorPmos: -1.40175e+08 muA
** NormalTransistorPmos: -8.30379e+07 muA
** NormalTransistorPmos: -1.40175e+08 muA
** NormalTransistorNmos: 8.30351e+07 muA
** NormalTransistorNmos: 8.30361e+07 muA
** NormalTransistorNmos: 8.30371e+07 muA
** NormalTransistorNmos: 8.30361e+07 muA
** NormalTransistorNmos: 1.14278e+08 muA
** DiodeTransistorNmos: 1.14277e+08 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 1.35721e+09 muA
** NormalTransistorNmos: 1.35721e+09 muA
** NormalTransistorPmos: -1.3572e+09 muA
** NormalTransistorPmos: -1.35721e+09 muA
** DiodeTransistorNmos: 1.19991e+07 muA
** NormalTransistorNmos: 1.19981e+07 muA
** DiodeTransistorNmos: 1.55771e+08 muA
** DiodeTransistorNmos: 1.58104e+08 muA
** DiodeTransistorPmos: -9.99589e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.10901  V
** inputVoltageBiasXXnXX3: 0.568001  V
** out: 2.5  V
** outFirstStage: 4.04001  V
** outInputVoltageBiasXXnXX1: 1.30201  V
** outSourceVoltageBiasXXnXX1: 0.652001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.704001  V
** innerTransistorStack1Load2: 0.525001  V
** innerTransistorStack2Load2: 0.525001  V
** sourceGCC1: 4.52501  V
** sourceGCC2: 4.52501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.363001  V
** innerTransconductance: 4.60401  V
** inner: 0.648001  V


.END