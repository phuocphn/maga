** Name: two_stage_single_output_op_amp_147_7

.MACRO two_stage_single_output_op_amp_147_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=12e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=407e-6
mSimpleFirstStageTransconductor5 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=14e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=66e-6
mSecondStage1StageBias8 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=12e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=14e-6
mMainBias11 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=168e-6
mSimpleFirstStageLoad12 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=294e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=358e-6
mSimpleFirstStageLoad14 outFirstStage outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=294e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12e-12
.EOM two_stage_single_output_op_amp_147_7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 5.11201 mW
** Area: 3237 (mu_m)^2
** Transit frequency: 5.16001 MHz
** Transit frequency with error factor: 5.14456 MHz
** Slew rate: 5.35819 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** VoutMax: 4.69001 V
** VoutMin: 0.150001 V
** VcmMax: 5.25 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 1.68134e+08 muA
** DiodeTransistorNmos: 8.95211e+07 muA
** DiodeTransistorNmos: 8.95221e+07 muA
** NormalTransistorNmos: 8.95211e+07 muA
** NormalTransistorNmos: 8.95221e+07 muA
** NormalTransistorPmos: -1.21893e+08 muA
** NormalTransistorPmos: -1.21893e+08 muA
** NormalTransistorNmos: 6.47451e+07 muA
** NormalTransistorNmos: 3.23721e+07 muA
** NormalTransistorNmos: 3.23721e+07 muA
** NormalTransistorNmos: 6.00477e+08 muA
** NormalTransistorPmos: -6.00476e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.68133e+08 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.12901  V
** outVoltageBiasXXpXX1: 4.28401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.09401  V
** innerTransistorStack2Load1: 1.09401  V
** sourceTransconductance: 1.92901  V


.END