** Name: two_stage_single_output_op_amp_161_4

.MACRO two_stage_single_output_op_amp_161_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=79e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=155e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=7e-6 W=259e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=24e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=255e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=255e-6
mSimpleFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=409e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=259e-6
mSecondStage1Transconductor10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=500e-6
mSimpleFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=409e-6
mSimpleFirstStageStageBias12 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=84e-6
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=129e-6
mSimpleFirstStageLoad14 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=7e-6 W=259e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=101e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=491e-6
mMainBias17 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=222e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=117e-6
mSecondStage1StageBias19 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=597e-6
mSimpleFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=7e-6 W=152e-6
mSimpleFirstStageTransconductor21 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=129e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.7001e-12
.EOM two_stage_single_output_op_amp_161_4

** Expected Performance Values: 
** Gain: 150 dB
** Power consumption: 6.25501 mW
** Area: 14694 (mu_m)^2
** Transit frequency: 3.72701 MHz
** Transit frequency with error factor: 3.72594 MHz
** Slew rate: 4.50159 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** VoutMax: 3.98001 V
** VoutMin: 0.370001 V
** VcmMax: 3.23001 V
** VcmMin: -0.25 V


** Expected Currents: 
** NormalTransistorPmos: -2.2508e+08 muA
** NormalTransistorPmos: -1.18622e+08 muA
** NormalTransistorPmos: -1.52165e+08 muA
** NormalTransistorPmos: -1.52165e+08 muA
** DiodeTransistorPmos: -1.52165e+08 muA
** NormalTransistorNmos: 1.94749e+08 muA
** NormalTransistorNmos: 1.94748e+08 muA
** NormalTransistorNmos: 1.94749e+08 muA
** NormalTransistorNmos: 1.94748e+08 muA
** NormalTransistorPmos: -8.51659e+07 muA
** NormalTransistorPmos: -8.51649e+07 muA
** NormalTransistorPmos: -4.25829e+07 muA
** NormalTransistorPmos: -4.25829e+07 muA
** NormalTransistorNmos: 4.97815e+08 muA
** NormalTransistorNmos: 4.97814e+08 muA
** NormalTransistorPmos: -4.97814e+08 muA
** NormalTransistorPmos: -4.97813e+08 muA
** DiodeTransistorNmos: 2.25081e+08 muA
** DiodeTransistorNmos: 1.18623e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.48201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.771001  V
** inputVoltageBiasXXnXX2: 0.569001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.26301  V
** innerTransistorStack1Load2: 0.216001  V
** innerTransistorStack2Load1: 3.95401  V
** innerTransistorStack2Load2: 0.216001  V
** out1: 2.76101  V
** sourceTransconductance: 3.25601  V
** innerStageBias: 4.26101  V
** innerTransconductance: 0.150001  V


.END