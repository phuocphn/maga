** Name: two_stage_single_output_op_amp_148_8

.MACRO two_stage_single_output_op_amp_148_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=10e-6 W=16e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias4 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=10e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=19e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=283e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=6e-6 W=570e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=10e-6 W=16e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=19e-6
mSimpleFirstStageLoad14 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=27e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=36e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=36e-6
mMainBias17 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=11e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=499e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=27e-6
mMainBias20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=30e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_148_8

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 4.07601 mW
** Area: 10795 (mu_m)^2
** Transit frequency: 2.51301 MHz
** Transit frequency with error factor: 2.51112 MHz
** Slew rate: 3.50005 V/mu_s
** Phase margin: 63.0254°
** CMRR: 109 dB
** VoutMax: 4.25 V
** VoutMin: 0.710001 V
** VcmMax: 4.54001 V
** VcmMin: 1.06001 V


** Expected Currents: 
** NormalTransistorPmos: -4.33469e+07 muA
** NormalTransistorPmos: -1.56479e+07 muA
** DiodeTransistorNmos: 4.35691e+07 muA
** DiodeTransistorNmos: 4.35691e+07 muA
** NormalTransistorNmos: 4.35681e+07 muA
** NormalTransistorNmos: 4.35691e+07 muA
** NormalTransistorPmos: -5.14729e+07 muA
** NormalTransistorPmos: -5.14729e+07 muA
** NormalTransistorPmos: -5.14719e+07 muA
** NormalTransistorPmos: -5.14729e+07 muA
** NormalTransistorNmos: 1.58071e+07 muA
** NormalTransistorNmos: 7.90301e+06 muA
** NormalTransistorNmos: 7.90301e+06 muA
** NormalTransistorNmos: 6.33318e+08 muA
** NormalTransistorNmos: 6.33317e+08 muA
** NormalTransistorPmos: -6.33317e+08 muA
** DiodeTransistorNmos: 4.33461e+07 muA
** DiodeTransistorNmos: 1.56471e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.835001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.03501  V
** outVoltageBiasXXnXX1: 1.11701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.10101  V
** innerTransistorStack1Load1: 1.12601  V
** innerTransistorStack1Load2: 4.15901  V
** innerTransistorStack2Load1: 1.12701  V
** innerTransistorStack2Load2: 4.15901  V
** sourceTransconductance: 1.87301  V
** innerStageBias: 0.430001  V


.END