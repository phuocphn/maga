** Name: two_stage_single_output_op_amp_71_7

.MACRO two_stage_single_output_op_amp_71_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=58e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=15e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=75e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=24e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=47e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=583e-6
mFoldedCascodeFirstStageLoad11 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=58e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=299e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=126e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=126e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=316e-6
mFoldedCascodeFirstStageLoad16 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=299e-6
mMainBias17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=130e-6
mMainBias18 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=423e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.40001e-12
.EOM two_stage_single_output_op_amp_71_7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 10.0661 mW
** Area: 6743 (mu_m)^2
** Transit frequency: 4.69401 MHz
** Transit frequency with error factor: 4.69041 MHz
** Slew rate: 5.39429 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** VoutMax: 4.25 V
** VoutMin: 0.180001 V
** VcmMax: 5.12001 V
** VcmMin: 1.5 V


** Expected Currents: 
** NormalTransistorPmos: -6.30879e+07 muA
** NormalTransistorPmos: -2.03663e+08 muA
** NormalTransistorPmos: -4.04779e+07 muA
** NormalTransistorPmos: -6.11469e+07 muA
** NormalTransistorPmos: -4.04779e+07 muA
** NormalTransistorPmos: -6.11469e+07 muA
** DiodeTransistorNmos: 4.04771e+07 muA
** NormalTransistorNmos: 4.04771e+07 muA
** NormalTransistorNmos: 4.13351e+07 muA
** NormalTransistorNmos: 4.13341e+07 muA
** NormalTransistorNmos: 2.06681e+07 muA
** NormalTransistorNmos: 2.06681e+07 muA
** NormalTransistorNmos: 1.60424e+09 muA
** NormalTransistorPmos: -1.60423e+09 muA
** DiodeTransistorNmos: 6.30871e+07 muA
** DiodeTransistorNmos: 2.03664e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** outVoltageBiasXXnXX1: 1.10701  V
** outVoltageBiasXXnXX2: 0.585001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.562001  V
** innerStageBias: 0.380001  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.90801  V


.END