** Name: two_stage_single_output_op_amp_147_11

.MACRO two_stage_single_output_op_amp_147_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=8e-6 W=18e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=31e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=14e-6
mMainBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=104e-6
mSecondStage1StageBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=25e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=177e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=33e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=31e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=55e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=201e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=18e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=33e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=120e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=337e-6
mSimpleFirstStageLoad16 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=90e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=220e-6
mMainBias18 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=386e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=600e-6
mSimpleFirstStageLoad20 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=90e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.20001e-12
.EOM two_stage_single_output_op_amp_147_11

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 7.60701 mW
** Area: 10988 (mu_m)^2
** Transit frequency: 3.40501 MHz
** Transit frequency with error factor: 3.38556 MHz
** Slew rate: 5.33456 V/mu_s
** Phase margin: 60.1606°
** CMRR: 87 dB
** VoutMax: 4.32001 V
** VoutMin: 0.540001 V
** VcmMax: 5.02001 V
** VcmMin: 0.840001 V


** Expected Currents: 
** NormalTransistorNmos: 8.46101e+07 muA
** NormalTransistorNmos: 2.39251e+08 muA
** NormalTransistorPmos: -5.18612e+08 muA
** DiodeTransistorNmos: 1.00399e+08 muA
** DiodeTransistorNmos: 1.004e+08 muA
** NormalTransistorNmos: 1.00399e+08 muA
** NormalTransistorNmos: 1.004e+08 muA
** NormalTransistorPmos: -1.19695e+08 muA
** NormalTransistorPmos: -1.19695e+08 muA
** NormalTransistorNmos: 3.85941e+07 muA
** NormalTransistorNmos: 1.92971e+07 muA
** NormalTransistorNmos: 1.92971e+07 muA
** NormalTransistorNmos: 4.29523e+08 muA
** NormalTransistorNmos: 4.29522e+08 muA
** NormalTransistorPmos: -4.29522e+08 muA
** NormalTransistorPmos: -4.29523e+08 muA
** DiodeTransistorNmos: 5.18613e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.46109e+07 muA
** DiodeTransistorPmos: -2.3925e+08 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.945001  V
** out: 2.5  V
** outFirstStage: 4.10401  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.04901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 0.961001  V
** innerTransistorStack2Load1: 0.961001  V
** sourceTransconductance: 1.84501  V
** innerStageBias: 0.183001  V
** innerTransconductance: 4.59501  V


.END