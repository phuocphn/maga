** Name: two_stage_single_output_op_amp_74_11

.MACRO two_stage_single_output_op_amp_74_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=39e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=8e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=12e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=36e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=323e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=39e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=46e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=46e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=36e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=574e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=12e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=9e-6 W=11e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=102e-6
mMainBias17 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=38e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=281e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=281e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=421e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=147e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=14e-6
mMainBias24 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=62e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_74_11

** Expected Performance Values: 
** Gain: 171 dB
** Power consumption: 3.96601 mW
** Area: 14985 (mu_m)^2
** Transit frequency: 5.15701 MHz
** Transit frequency with error factor: 5.15718 MHz
** Slew rate: 4.86045 V/mu_s
** Phase margin: 69.9009°
** CMRR: 133 dB
** VoutMax: 4.26001 V
** VoutMin: 0.710001 V
** VcmMax: 5.15001 V
** VcmMin: 1.47001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorNmos: 3.72781e+07 muA
** NormalTransistorPmos: -7.24799e+06 muA
** NormalTransistorPmos: -2.19049e+07 muA
** NormalTransistorPmos: -3.28559e+07 muA
** NormalTransistorPmos: -2.19079e+07 muA
** NormalTransistorPmos: -3.28609e+07 muA
** NormalTransistorNmos: 2.19061e+07 muA
** NormalTransistorNmos: 2.19071e+07 muA
** DiodeTransistorNmos: 2.19061e+07 muA
** NormalTransistorNmos: 2.19031e+07 muA
** DiodeTransistorNmos: 2.19021e+07 muA
** NormalTransistorNmos: 1.09521e+07 muA
** NormalTransistorNmos: 1.09521e+07 muA
** NormalTransistorNmos: 5.71389e+08 muA
** NormalTransistorNmos: 5.71388e+08 muA
** NormalTransistorPmos: -5.71388e+08 muA
** NormalTransistorPmos: -5.71389e+08 muA
** DiodeTransistorNmos: 7.24701e+06 muA
** NormalTransistorNmos: 7.24601e+06 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -3.72789e+07 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.16001  V
** outInputVoltageBiasXXnXX1: 1.31801  V
** outSourceVoltageBiasXXnXX1: 0.659001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.18101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.620001  V
** out1: 1.48301  V
** sourceGCC1: 4.54501  V
** sourceGCC2: 4.54501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.579001  V
** innerTransconductance: 4.71501  V
** inner: 0.659001  V


.END