** Name: two_stage_single_output_op_amp_80_1

.MACRO two_stage_single_output_op_amp_80_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=12e-6
mFoldedCascodeFirstStageStageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=172e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=74e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=49e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=45e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=163e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=163e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=99e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=99e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=172e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mSecondStage1Transconductor13 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=348e-6
mFoldedCascodeFirstStageLoad14 outFirstStage outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=45e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=455e-6
mMainBias16 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=140e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=329e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=74e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=74e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=595e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=329e-6
mMainBias22 outVoltageBiasXXnXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=195e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.8001e-12
.EOM two_stage_single_output_op_amp_80_1

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 13.5631 mW
** Area: 8681 (mu_m)^2
** Transit frequency: 7.11501 MHz
** Transit frequency with error factor: 7.11526 MHz
** Slew rate: 5.25327 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.64001 V
** VoutMin: 0.310001 V
** VcmMax: 5.04001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 3.75676e+08 muA
** NormalTransistorNmos: 1.15905e+08 muA
** NormalTransistorPmos: -4.53561e+08 muA
** NormalTransistorPmos: -1.04397e+08 muA
** NormalTransistorPmos: -1.75039e+08 muA
** NormalTransistorPmos: -1.04397e+08 muA
** NormalTransistorPmos: -1.75039e+08 muA
** NormalTransistorNmos: 1.04398e+08 muA
** NormalTransistorNmos: 1.04397e+08 muA
** NormalTransistorNmos: 1.04398e+08 muA
** NormalTransistorNmos: 1.04397e+08 muA
** NormalTransistorNmos: 1.41288e+08 muA
** DiodeTransistorNmos: 1.41289e+08 muA
** NormalTransistorNmos: 7.06431e+07 muA
** NormalTransistorNmos: 7.06431e+07 muA
** NormalTransistorNmos: 1.40742e+09 muA
** NormalTransistorPmos: -1.40741e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 4.53562e+08 muA
** DiodeTransistorPmos: -3.75675e+08 muA
** DiodeTransistorPmos: -1.15904e+08 muA


** Expected Voltages: 
** ibias: 1.20501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.715001  V
** outSourceVoltageBiasXXnXX1: 0.603001  V
** outVoltageBiasXXnXX2: 0.920001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.07401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 4.43801  V
** sourceGCC2: 4.43801  V
** sourceTransconductance: 1.93601  V
** inner: 0.601001  V


.END