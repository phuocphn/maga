** Name: two_stage_single_output_op_amp_162_4

.MACRO two_stage_single_output_op_amp_162_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=47e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=5e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=4e-6 W=53e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=157e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=240e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=93e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=93e-6
mSimpleFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=5e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=597e-6
mSecondStage1Transconductor12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=35e-6
mSimpleFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=5e-6
mMainBias14 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=79e-6
mSimpleFirstStageTransconductor15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=21e-6
mSimpleFirstStageLoad16 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=5e-6
mSimpleFirstStageStageBias17 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=240e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=64e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=157e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSecondStage1StageBias21 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=4e-6 W=600e-6
mSimpleFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=11e-6
mSimpleFirstStageTransconductor23 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=21e-6
mMainBias24 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=23e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_162_4

** Expected Performance Values: 
** Gain: 145 dB
** Power consumption: 1.53601 mW
** Area: 14990 (mu_m)^2
** Transit frequency: 3.46401 MHz
** Transit frequency with error factor: 3.46065 MHz
** Slew rate: 5.69031 V/mu_s
** Phase margin: 62.4525°
** CMRR: 94 dB
** VoutMax: 3.44001 V
** VoutMin: 0.480001 V
** VcmMax: 3.23001 V
** VcmMin: -0.109999 V


** Expected Currents: 
** NormalTransistorNmos: 1.67191e+07 muA
** NormalTransistorPmos: -5.83819e+07 muA
** NormalTransistorPmos: -9.95299e+06 muA
** NormalTransistorPmos: -7.05599e+06 muA
** NormalTransistorPmos: -7.05599e+06 muA
** DiodeTransistorPmos: -7.05599e+06 muA
** NormalTransistorNmos: 1.98801e+07 muA
** NormalTransistorNmos: 1.98791e+07 muA
** NormalTransistorNmos: 1.98801e+07 muA
** NormalTransistorNmos: 1.98791e+07 muA
** NormalTransistorPmos: -2.56509e+07 muA
** DiodeTransistorPmos: -2.56519e+07 muA
** NormalTransistorPmos: -1.28249e+07 muA
** NormalTransistorPmos: -1.28249e+07 muA
** NormalTransistorNmos: 1.62455e+08 muA
** NormalTransistorNmos: 1.62454e+08 muA
** NormalTransistorPmos: -1.62454e+08 muA
** NormalTransistorPmos: -1.62453e+08 muA
** DiodeTransistorNmos: 5.83811e+07 muA
** DiodeTransistorNmos: 9.95201e+06 muA
** DiodeTransistorPmos: -1.67199e+07 muA
** NormalTransistorPmos: -1.67209e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.91601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.49201  V
** outSourceVoltageBiasXXpXX1: 4.24601  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX1: 0.885001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.80501  V
** innerTransistorStack1Load2: 0.172001  V
** innerTransistorStack2Load2: 0.172001  V
** out1: 3.05101  V
** sourceTransconductance: 3.32501  V
** innerStageBias: 3.72501  V
** innerTransconductance: 0.150001  V
** inner: 4.24501  V


.END