** Name: symmetrical_op_amp114

.MACRO symmetrical_op_amp114 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias4 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=257e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=6e-6 W=24e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mSymmetricalFirstStageTransconductor8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=15e-6
mSecondStage1StageBias9 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=34e-6
mSymmetricalFirstStageTransconductor10 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=15e-6
mMainBias11 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=6e-6 W=18e-6
mMainBias12 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=59e-6
mSymmetricalFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=13e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=13e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=35e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=35e-6
mSymmetricalFirstStageLoad17 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=83e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=224e-6
mSecondStage1Transconductor19 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=224e-6
mSymmetricalFirstStageLoad20 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=83e-6
mMainBias21 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=363e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp114

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 1.78801 mW
** Area: 3836 (mu_m)^2
** Transit frequency: 3.125 MHz
** Transit frequency with error factor: 3.12456 MHz
** Slew rate: 4.53596 V/mu_s
** Phase margin: 80.7871°
** CMRR: 140 dB
** negPSRR: 134 dB
** posPSRR: 62 dB
** VoutMax: 4.25 V
** VoutMin: 0.360001 V
** VcmMax: 4.81001 V
** VcmMin: 0.950001 V


** Expected Currents: 
** NormalTransistorNmos: 8.28191e+07 muA
** NormalTransistorNmos: 2.53821e+07 muA
** NormalTransistorPmos: -1.1483e+08 muA
** NormalTransistorPmos: -1.68449e+07 muA
** NormalTransistorPmos: -1.68459e+07 muA
** NormalTransistorPmos: -1.68449e+07 muA
** NormalTransistorPmos: -1.68459e+07 muA
** NormalTransistorNmos: 3.36891e+07 muA
** NormalTransistorNmos: 1.68441e+07 muA
** NormalTransistorNmos: 1.68441e+07 muA
** NormalTransistorNmos: 4.54861e+07 muA
** NormalTransistorNmos: 4.54851e+07 muA
** NormalTransistorPmos: -4.54869e+07 muA
** NormalTransistorPmos: -4.54869e+07 muA
** DiodeTransistorNmos: 4.54861e+07 muA
** NormalTransistorPmos: -4.54869e+07 muA
** NormalTransistorPmos: -4.54869e+07 muA
** DiodeTransistorNmos: 1.14831e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.28199e+07 muA
** DiodeTransistorPmos: -2.53829e+07 muA


** Expected Voltages: 
** ibias: 0.722001  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.588001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 1.13801  V
** outVoltageBiasXXpXX0: 4.24701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.86401  V
** innerStageBias: 0.555001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END