** Name: one_stage_single_output_op_amp79

.MACRO one_stage_single_output_op_amp79 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=36e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageStageBias5 FirstStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=54e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=46e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=46e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=57e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=83e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=83e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=97e-6
mFoldedCascodeFirstStageLoad12 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=57e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=111e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=111e-6
mMainBias16 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mFoldedCascodeFirstStageLoad17 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=600e-6
mMainBias18 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=129e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp79

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 3.84801 mW
** Area: 4596 (mu_m)^2
** Transit frequency: 5.20001 MHz
** Transit frequency with error factor: 5.19994 MHz
** Slew rate: 6.62351 V/mu_s
** Phase margin: 83.6519°
** CMRR: 140 dB
** VoutMax: 3.80001 V
** VoutMin: 0.350001 V
** VcmMax: 4.93001 V
** VcmMin: 1.44001 V


** Expected Currents: 
** NormalTransistorPmos: -2.59594e+08 muA
** NormalTransistorPmos: -3.8e+07 muA
** NormalTransistorPmos: -1.33477e+08 muA
** NormalTransistorPmos: -2.2603e+08 muA
** NormalTransistorPmos: -1.33477e+08 muA
** NormalTransistorPmos: -2.2603e+08 muA
** NormalTransistorNmos: 1.33478e+08 muA
** NormalTransistorNmos: 1.33477e+08 muA
** NormalTransistorNmos: 1.33478e+08 muA
** NormalTransistorNmos: 1.33477e+08 muA
** NormalTransistorNmos: 1.85104e+08 muA
** NormalTransistorNmos: 1.85103e+08 muA
** NormalTransistorNmos: 9.25521e+07 muA
** NormalTransistorNmos: 9.25521e+07 muA
** DiodeTransistorNmos: 2.59595e+08 muA
** DiodeTransistorNmos: 3.79991e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.22001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.606001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 3.96101  V
** outVoltageBiasXXnXX1: 0.956001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.401001  V
** innerTransistorStack1Load2: 0.384001  V
** innerTransistorStack2Load2: 0.385001  V
** out1: 0.590001  V
** sourceGCC1: 3.94101  V
** sourceGCC2: 3.94101  V
** sourceTransconductance: 1.81301  V


.END