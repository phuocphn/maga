** Name: two_stage_single_output_op_amp_29_11

.MACRO two_stage_single_output_op_amp_29_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=7e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=523e-6
mSecondStage1StageBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
mSimpleFirstStageStageBias5 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=313e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=29e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=225e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=400e-6
mSecondStage1StageBias9 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=300e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=29e-6
mMainBias11 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=422e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=599e-6
mSecondStage1Transconductor13 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=523e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.6001e-12
.EOM two_stage_single_output_op_amp_29_11

** Expected Performance Values: 
** Gain: 132 dB
** Power consumption: 5.64601 mW
** Area: 7208 (mu_m)^2
** Transit frequency: 6.08301 MHz
** Transit frequency with error factor: 6.04811 MHz
** Slew rate: 12.7761 V/mu_s
** Phase margin: 60.1606°
** CMRR: 87 dB
** negPSRR: 113 dB
** posPSRR: 85 dB
** VoutMax: 4.62001 V
** VoutMin: 0.730001 V
** VcmMax: 4.66001 V
** VcmMin: 1.89001 V


** Expected Currents: 
** NormalTransistorNmos: 4.16289e+08 muA
** DiodeTransistorPmos: -1.54678e+08 muA
** NormalTransistorPmos: -1.54678e+08 muA
** NormalTransistorNmos: 3.09356e+08 muA
** NormalTransistorNmos: 3.09355e+08 muA
** NormalTransistorNmos: 1.54679e+08 muA
** NormalTransistorNmos: 1.54679e+08 muA
** NormalTransistorNmos: 3.93492e+08 muA
** NormalTransistorNmos: 3.93491e+08 muA
** NormalTransistorPmos: -3.93491e+08 muA
** NormalTransistorPmos: -3.93492e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -4.16288e+08 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.24401  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.560001  V
** out1: 4.25401  V
** sourceTransconductance: 1.34501  V
** innerStageBias: 0.565001  V
** innerTransconductance: 4.44101  V


.END