** Name: one_stage_single_output_op_amp119

.MACRO one_stage_single_output_op_amp119 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=6e-6
mMainBias2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=15e-6
mTelescopicFirstStageLoad4 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=58e-6
mTelescopicFirstStageLoad5 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=43e-6
mTelescopicFirstStageLoad7 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=111e-6
mTelescopicFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=78e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=16e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=16e-6
mTelescopicFirstStageLoad11 out outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=111e-6
mMainBias12 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mTelescopicFirstStageStageBias13 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=81e-6
mTelescopicFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad15 out FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=58e-6
mMainBias16 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=89e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp119

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 0.475001 mW
** Area: 2853 (mu_m)^2
** Transit frequency: 3.22401 MHz
** Transit frequency with error factor: 3.22421 MHz
** Slew rate: 3.84589 V/mu_s
** Phase margin: 80.7871°
** CMRR: 153 dB
** VoutMax: 3.85001 V
** VoutMin: 0.600001 V
** VcmMax: 3.54001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 7.92701e+06 muA
** NormalTransistorPmos: -1.61879e+07 muA
** NormalTransistorNmos: 3.04741e+07 muA
** NormalTransistorNmos: 3.04741e+07 muA
** DiodeTransistorPmos: -3.04749e+07 muA
** DiodeTransistorPmos: -3.04759e+07 muA
** NormalTransistorPmos: -3.04749e+07 muA
** NormalTransistorPmos: -3.04759e+07 muA
** NormalTransistorNmos: 7.71381e+07 muA
** NormalTransistorNmos: 7.71371e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** DiodeTransistorNmos: 1.61871e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.92799e+06 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 4.21001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerOutputLoad2: 3.28501  V
** innerStageBias: 0.606001  V
** innerTransistorStack1Load2: 4.02101  V
** innerTransistorStack2Load2: 4.02001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END