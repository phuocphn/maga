** Name: two_stage_single_output_op_amp_24_6

.MACRO two_stage_single_output_op_amp_24_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias3 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=7e-6 W=20e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=531e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=129e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=354e-6
mSimpleFirstStageLoad7 FirstStageYinnerSourceLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=36e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=129e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=129e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=375e-6
mSecondStage1Transconductor11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=98e-6
mSimpleFirstStageLoad12 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=36e-6
mMainBias13 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=77e-6
mSimpleFirstStageTransconductor14 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=51e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=129e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=531e-6
mMainBias17 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=20e-6
mSecondStage1StageBias18 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=7e-6 W=354e-6
mSimpleFirstStageTransconductor19 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=51e-6
mMainBias20 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=70e-6
mMainBias21 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=36e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_24_6

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 2.67901 mW
** Area: 12241 (mu_m)^2
** Transit frequency: 4.96301 MHz
** Transit frequency with error factor: 4.95393 MHz
** Slew rate: 7.31431 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** negPSRR: 95 dB
** posPSRR: 103 dB
** VoutMax: 3.54001 V
** VoutMin: 0.400001 V
** VcmMax: 3.18001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.27312e+08 muA
** NormalTransistorPmos: -3.55839e+07 muA
** NormalTransistorPmos: -1.82999e+07 muA
** NormalTransistorNmos: 2.72991e+07 muA
** NormalTransistorNmos: 2.73001e+07 muA
** NormalTransistorNmos: 2.72991e+07 muA
** NormalTransistorNmos: 2.73001e+07 muA
** NormalTransistorPmos: -5.46009e+07 muA
** DiodeTransistorPmos: -5.46019e+07 muA
** NormalTransistorPmos: -2.72999e+07 muA
** NormalTransistorPmos: -2.72999e+07 muA
** NormalTransistorNmos: 1.79954e+08 muA
** NormalTransistorNmos: 1.79953e+08 muA
** NormalTransistorPmos: -1.79953e+08 muA
** DiodeTransistorPmos: -1.79952e+08 muA
** DiodeTransistorNmos: 3.55831e+07 muA
** DiodeTransistorNmos: 1.82991e+07 muA
** DiodeTransistorPmos: -2.27311e+08 muA
** NormalTransistorPmos: -2.27312e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.98001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.56401  V
** outSourceVoltageBiasXXpXX1: 4.28201  V
** outSourceVoltageBiasXXpXX2: 3.99201  V
** outVoltageBiasXXnXX0: 0.592001  V
** outVoltageBiasXXnXX1: 0.809001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.240001  V
** innerTransistorStack2Load1: 0.240001  V
** sourceTransconductance: 3.45001  V
** innerTransconductance: 0.150001  V
** inner: 4.28201  V
** inner: 3.98501  V


.END