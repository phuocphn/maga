** Name: symmetrical_op_amp37

.MACRO symmetrical_op_amp37 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=111e-6
mMainBias6 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=34e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=34e-6
mMainBias9 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=52e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=20e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=20e-6
mSymmetricalFirstStageStageBias12 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=245e-6
mSymmetricalFirstStageStageBias13 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=52e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias15 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mMainBias16 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=7e-6 W=354e-6
mSymmetricalFirstStageTransconductor17 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=49e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias18 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=1e-6 W=17e-6
mMainBias19 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=210e-6
mSecondStage1StageBias20 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageTransconductor21 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=49e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp37

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 1.31301 mW
** Area: 7517 (mu_m)^2
** Transit frequency: 3.43701 MHz
** Transit frequency with error factor: 3.43673 MHz
** Slew rate: 3.50006 V/mu_s
** Phase margin: 77.3494°
** CMRR: 143 dB
** negPSRR: 50 dB
** posPSRR: 57 dB
** VoutMax: 4.35001 V
** VoutMin: 0.570001 V
** VcmMax: 3.37001 V
** VcmMin: 0.0600001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00041e+08 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -3.18819e+07 muA
** DiodeTransistorNmos: 1.11561e+07 muA
** DiodeTransistorNmos: 1.11541e+07 muA
** NormalTransistorPmos: -2.23109e+07 muA
** NormalTransistorPmos: -2.23119e+07 muA
** NormalTransistorPmos: -1.11549e+07 muA
** NormalTransistorPmos: -1.11549e+07 muA
** NormalTransistorNmos: 3.50111e+07 muA
** NormalTransistorNmos: 3.50101e+07 muA
** NormalTransistorPmos: -3.50119e+07 muA
** NormalTransistorPmos: -3.50129e+07 muA
** NormalTransistorPmos: -3.43309e+07 muA
** NormalTransistorPmos: -3.43319e+07 muA
** NormalTransistorNmos: 3.43301e+07 muA
** NormalTransistorNmos: 3.43291e+07 muA
** DiodeTransistorNmos: 1.90471e+07 muA
** DiodeTransistorNmos: 3.18811e+07 muA
** DiodeTransistorPmos: -1.0004e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24801  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 3.68601  V
** inOutputTransconductanceComplementarySecondStage: 0.976001  V
** inSourceTransconductanceComplementarySecondStage: 0.624001  V
** innerComplementarySecondStage: 4.22601  V
** inputVoltageBiasXXnXX0: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.625  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40501  V
** sourceTransconductance: 3.22301  V
** innerStageBias: 4.69101  V
** innerTransconductance: 0.220001  V
** inner: 4.58501  V
** inner: 0.221001  V


.END