** Name: two_stage_single_output_op_amp_10_7

.MACRO two_stage_single_output_op_amp_10_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=13e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mSimpleFirstStageTransconductor4 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=9e-6
mSimpleFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mMainBias6 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=54e-6
mSecondStage1StageBias7 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=343e-6
mSimpleFirstStageTransconductor8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=9e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=13e-6
mSecondStage1Transconductor10 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=297e-6
mSimpleFirstStageLoad11 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=59e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_10_7

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 2.96201 mW
** Area: 2468 (mu_m)^2
** Transit frequency: 2.74101 MHz
** Transit frequency with error factor: 2.73858 MHz
** Slew rate: 5.27925 V/mu_s
** Phase margin: 68.182°
** CMRR: 92 dB
** negPSRR: 136 dB
** posPSRR: 90 dB
** VoutMax: 4.40001 V
** VoutMin: 0.180001 V
** VcmMax: 4.09001 V
** VcmMin: 0.900001 V


** Expected Currents: 
** NormalTransistorNmos: 7.61491e+07 muA
** DiodeTransistorPmos: -1.19299e+07 muA
** NormalTransistorPmos: -1.19299e+07 muA
** NormalTransistorPmos: -1.19299e+07 muA
** NormalTransistorNmos: 2.38581e+07 muA
** NormalTransistorNmos: 1.19291e+07 muA
** NormalTransistorNmos: 1.19291e+07 muA
** NormalTransistorNmos: 4.82489e+08 muA
** NormalTransistorPmos: -4.82488e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.61499e+07 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.83601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.83601  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.78701  V


.END