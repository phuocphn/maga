** Name: two_stage_single_output_op_amp_187_12

.MACRO two_stage_single_output_op_amp_187_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=8e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=29e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=372e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSecondStage1StageBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=237e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=178e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=187e-6
mSimpleFirstStageLoad10 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=50e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=29e-6
mMainBias13 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=262e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=372e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=13e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=187e-6
mMainBias17 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=151e-6
mSimpleFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=576e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=559e-6
mSecondStage1Transconductor20 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad21 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=576e-6
mMainBias22 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=272e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.7001e-12
.EOM two_stage_single_output_op_amp_187_12

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 11.6971 mW
** Area: 13364 (mu_m)^2
** Transit frequency: 9.06501 MHz
** Transit frequency with error factor: 9.04108 MHz
** Slew rate: 8.54367 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 0.830001 V
** VcmMax: 5.10001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 1.72607e+08 muA
** NormalTransistorNmos: 9.94881e+07 muA
** NormalTransistorPmos: -1.14181e+08 muA
** NormalTransistorNmos: 1.78867e+08 muA
** NormalTransistorNmos: 1.78868e+08 muA
** DiodeTransistorNmos: 1.78867e+08 muA
** NormalTransistorPmos: -2.38227e+08 muA
** NormalTransistorPmos: -2.38227e+08 muA
** NormalTransistorNmos: 1.18722e+08 muA
** NormalTransistorNmos: 1.18721e+08 muA
** NormalTransistorNmos: 5.93611e+07 muA
** NormalTransistorNmos: 5.93611e+07 muA
** NormalTransistorNmos: 1.46669e+09 muA
** DiodeTransistorNmos: 1.46669e+09 muA
** NormalTransistorPmos: -1.46668e+09 muA
** NormalTransistorPmos: -1.46668e+09 muA
** DiodeTransistorNmos: 1.14182e+08 muA
** NormalTransistorNmos: 1.14181e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.72606e+08 muA
** DiodeTransistorPmos: -9.94889e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.05401  V
** outInputVoltageBiasXXnXX1: 1.24001  V
** outSourceVoltageBiasXXnXX1: 0.620001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX2: 4.13101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.477001  V
** innerTransistorStack2Load1: 1.15501  V
** out1: 2.13301  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.61801  V
** inner: 0.619001  V


.END