** Name: symmetrical_op_amp116

.MACRO symmetrical_op_amp116 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=11e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias3 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=9e-6
mSymmetricalFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=96e-6
mSecondStage1StageBias6 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=45e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias7 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=45e-6
mSymmetricalFirstStageTransconductor8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=47e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias9 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=2e-6 W=91e-6
mSecondStage1StageBias10 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=91e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=47e-6
mMainBias12 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=7e-6 W=28e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=16e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mSymmetricalFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=43e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=43e-6
mMainBias18 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=19e-6
mSymmetricalFirstStageLoad19 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=211e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor20 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=463e-6
mSecondStage1Transconductor21 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=463e-6
mSymmetricalFirstStageLoad22 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=211e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp116

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 1.75601 mW
** Area: 5239 (mu_m)^2
** Transit frequency: 7.02101 MHz
** Transit frequency with error factor: 7.02112 MHz
** Slew rate: 9.25896 V/mu_s
** Phase margin: 77.3494°
** CMRR: 142 dB
** negPSRR: 111 dB
** posPSRR: 62 dB
** VoutMax: 4.25 V
** VoutMin: 0.380001 V
** VcmMax: 4.81001 V
** VcmMin: 0.890001 V


** Expected Currents: 
** NormalTransistorNmos: 1.43091e+07 muA
** NormalTransistorNmos: 2.53821e+07 muA
** NormalTransistorPmos: -2.96239e+07 muA
** NormalTransistorPmos: -4.28339e+07 muA
** NormalTransistorPmos: -4.28349e+07 muA
** NormalTransistorPmos: -4.28339e+07 muA
** NormalTransistorPmos: -4.28349e+07 muA
** NormalTransistorNmos: 8.56661e+07 muA
** NormalTransistorNmos: 4.28331e+07 muA
** NormalTransistorNmos: 4.28331e+07 muA
** NormalTransistorNmos: 9.31401e+07 muA
** NormalTransistorNmos: 9.31391e+07 muA
** NormalTransistorPmos: -9.31409e+07 muA
** NormalTransistorPmos: -9.31399e+07 muA
** NormalTransistorNmos: 9.31401e+07 muA
** NormalTransistorNmos: 9.31391e+07 muA
** NormalTransistorPmos: -9.31409e+07 muA
** NormalTransistorPmos: -9.31399e+07 muA
** DiodeTransistorNmos: 2.96231e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.43099e+07 muA
** DiodeTransistorPmos: -2.53829e+07 muA


** Expected Voltages: 
** ibias: 0.678001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.781001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.626001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 3.70901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.88701  V
** innerStageBias: 0.221001  V
** innerTransconductance: 4.40001  V
** inner: 0.221001  V
** inner: 4.40001  V


.END