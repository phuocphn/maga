** Name: two_stage_single_output_op_amp_152_11

.MACRO two_stage_single_output_op_amp_152_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=24e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=113e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=46e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=511e-6
mMainBias11 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=14e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=563e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=24e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=113e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=87e-6
mSimpleFirstStageLoad16 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=214e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=472e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=472e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=424e-6
mMainBias20 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=146e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=214e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.5e-12
.EOM two_stage_single_output_op_amp_152_11

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 14.8921 mW
** Area: 9215 (mu_m)^2
** Transit frequency: 7.49501 MHz
** Transit frequency with error factor: 7.4908 MHz
** Slew rate: 7.23022 V/mu_s
** Phase margin: 60.1606°
** CMRR: 118 dB
** VoutMax: 4.25 V
** VoutMin: 0.710001 V
** VcmMax: 4.73001 V
** VcmMin: 0.900001 V


** Expected Currents: 
** NormalTransistorNmos: 2.13221e+08 muA
** NormalTransistorNmos: 3.50031e+07 muA
** NormalTransistorPmos: -1.96602e+08 muA
** DiodeTransistorNmos: 5.75737e+08 muA
** NormalTransistorNmos: 5.75738e+08 muA
** NormalTransistorNmos: 5.75739e+08 muA
** DiodeTransistorNmos: 5.75738e+08 muA
** NormalTransistorPmos: -6.32103e+08 muA
** NormalTransistorPmos: -6.32104e+08 muA
** NormalTransistorPmos: -6.32105e+08 muA
** NormalTransistorPmos: -6.32104e+08 muA
** NormalTransistorNmos: 1.12736e+08 muA
** NormalTransistorNmos: 5.63671e+07 muA
** NormalTransistorNmos: 5.63671e+07 muA
** NormalTransistorNmos: 1.25936e+09 muA
** NormalTransistorNmos: 1.25936e+09 muA
** NormalTransistorPmos: -1.25935e+09 muA
** NormalTransistorPmos: -1.25935e+09 muA
** DiodeTransistorNmos: 1.96603e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.1322e+08 muA
** DiodeTransistorPmos: -3.50039e+07 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11201  V
** inputVoltageBiasXXpXX2: 4.16101  V
** out: 2.5  V
** outFirstStage: 4.02701  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerTransistorStack1Load1: 1.15601  V
** innerTransistorStack1Load2: 4.65501  V
** innerTransistorStack2Load1: 1.15501  V
** innerTransistorStack2Load2: 4.65501  V
** sourceTransconductance: 1.94101  V
** innerStageBias: 0.342001  V
** innerTransconductance: 4.59101  V


.END