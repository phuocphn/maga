** Name: two_stage_single_output_op_amp_72_8

.MACRO two_stage_single_output_op_amp_72_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=22e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=60e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=20e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=39e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=13e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=30e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=30e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=39e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=184e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=60e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=7e-6 W=143e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=22e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=51e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=593e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=51e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=35e-6
mMainBias21 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=61e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_72_8

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 5.20601 mW
** Area: 8221 (mu_m)^2
** Transit frequency: 4.99401 MHz
** Transit frequency with error factor: 4.98884 MHz
** Slew rate: 4.21016 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** VoutMax: 4.25 V
** VoutMin: 1.73001 V
** VcmMax: 5.17001 V
** VcmMin: 1.30001 V


** Expected Currents: 
** NormalTransistorPmos: -3.54849e+07 muA
** NormalTransistorPmos: -6.06219e+07 muA
** NormalTransistorPmos: -2.07119e+07 muA
** NormalTransistorPmos: -3.24439e+07 muA
** NormalTransistorPmos: -2.07119e+07 muA
** NormalTransistorPmos: -3.24439e+07 muA
** DiodeTransistorNmos: 2.07111e+07 muA
** NormalTransistorNmos: 2.07111e+07 muA
** NormalTransistorNmos: 2.34611e+07 muA
** DiodeTransistorNmos: 2.34601e+07 muA
** NormalTransistorNmos: 1.17311e+07 muA
** NormalTransistorNmos: 1.17311e+07 muA
** NormalTransistorNmos: 8.60138e+08 muA
** NormalTransistorNmos: 8.60137e+08 muA
** NormalTransistorPmos: -8.60137e+08 muA
** DiodeTransistorNmos: 3.54841e+07 muA
** NormalTransistorNmos: 3.54831e+07 muA
** DiodeTransistorNmos: 6.06211e+07 muA
** DiodeTransistorNmos: 6.06201e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.14601  V
** outInputVoltageBiasXXnXX2: 1.92801  V
** outSourceVoltageBiasXXnXX1: 0.573001  V
** outSourceVoltageBiasXXnXX2: 1.02401  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.615001  V
** sourceGCC1: 4.11201  V
** sourceGCC2: 4.11201  V
** sourceTransconductance: 1.94301  V
** innerStageBias: 0.819001  V
** inner: 0.573001  V


.END