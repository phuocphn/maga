** Name: two_stage_single_output_op_amp_54_9

.MACRO two_stage_single_output_op_amp_54_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=24e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=69e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=401e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=19e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=26e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=14e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=119e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=119e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=25e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=25e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=401e-6
mFoldedCascodeFirstStageLoad15 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=14e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=169e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=88e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=88e-6
mMainBias19 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=200e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=327e-6
mMainBias21 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=365e-6
mSecondStage1Transconductor22 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=254e-6
mFoldedCascodeFirstStageLoad23 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=169e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_54_9

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 8.60401 mW
** Area: 8547 (mu_m)^2
** Transit frequency: 4.42801 MHz
** Transit frequency with error factor: 4.42829 MHz
** Slew rate: 4.99915 V/mu_s
** Phase margin: 61.8795°
** CMRR: 147 dB
** VoutMax: 4.25 V
** VoutMin: 0.790001 V
** VcmMax: 5.15001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorPmos: -7.72349e+07 muA
** NormalTransistorPmos: -1.24929e+08 muA
** NormalTransistorPmos: -1.40736e+08 muA
** NormalTransistorPmos: -2.27739e+07 muA
** NormalTransistorPmos: -3.41599e+07 muA
** NormalTransistorPmos: -2.27739e+07 muA
** NormalTransistorPmos: -3.41599e+07 muA
** NormalTransistorNmos: 2.27731e+07 muA
** NormalTransistorNmos: 2.27721e+07 muA
** NormalTransistorNmos: 2.27731e+07 muA
** NormalTransistorNmos: 2.27721e+07 muA
** NormalTransistorNmos: 2.27731e+07 muA
** NormalTransistorNmos: 1.13871e+07 muA
** NormalTransistorNmos: 1.13871e+07 muA
** NormalTransistorNmos: 1.28949e+09 muA
** DiodeTransistorNmos: 1.28949e+09 muA
** NormalTransistorPmos: -1.28948e+09 muA
** DiodeTransistorNmos: 7.72341e+07 muA
** NormalTransistorNmos: 7.72331e+07 muA
** DiodeTransistorNmos: 1.2493e+08 muA
** DiodeTransistorNmos: 1.40737e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.19801  V
** inputVoltageBiasXXnXX2: 0.951001  V
** inputVoltageBiasXXnXX3: 0.561001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.599001  V
** outSourceVoltageBiasXXpXX1: 4.18201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.91501  V
** inner: 0.598001  V


.END