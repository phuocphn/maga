** Name: symmetrical_op_amp147

.MACRO symmetrical_op_amp147 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias3 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=104e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=3e-6 W=104e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=159e-6
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=159e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=154e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=154e-6
mSymmetricalFirstStageLoad10 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=70e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=1e-6 W=68e-6
mSecondStage1Transconductor12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=68e-6
mSymmetricalFirstStageLoad13 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=70e-6
mSymmetricalFirstStageStageBias14 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSymmetricalFirstStageStageBias15 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=518e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias16 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=104e-6
mSymmetricalFirstStageTransconductor17 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=420e-6
mSecondStage1StageBias18 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=3e-6 W=104e-6
mSymmetricalFirstStageTransconductor19 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=420e-6
mMainBias20 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=193e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp147

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 7.05301 mW
** Area: 5177 (mu_m)^2
** Transit frequency: 16.4361 MHz
** Transit frequency with error factor: 16.436 MHz
** Slew rate: 29.488 V/mu_s
** Phase margin: 85.3708°
** CMRR: 139 dB
** negPSRR: 46 dB
** posPSRR: 167 dB
** VoutMax: 3.05001 V
** VoutMin: 0.380001 V
** VcmMax: 3.10001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.93413e+08 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04163e+08 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04163e+08 muA
** NormalTransistorPmos: -6.08327e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorNmos: 2.95474e+08 muA
** NormalTransistorNmos: 2.95473e+08 muA
** NormalTransistorPmos: -2.95473e+08 muA
** DiodeTransistorPmos: -2.95474e+08 muA
** DiodeTransistorPmos: -2.93312e+08 muA
** NormalTransistorPmos: -2.93313e+08 muA
** NormalTransistorNmos: 2.93313e+08 muA
** NormalTransistorNmos: 2.93314e+08 muA
** DiodeTransistorNmos: 1.93414e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 3.74501  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 2.48701  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.781001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.21801  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.34801  V
** innerTransconductance: 0.150001  V
** inner: 3.73601  V
** inner: 0.150001  V


.END