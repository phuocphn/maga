** Name: symmetrical_op_amp149

.MACRO symmetrical_op_amp149 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=15e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=34e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=70e-6
mSymmetricalFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=317e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=5e-6
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=124e-6
mSymmetricalFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=123e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=114e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=114e-6
mSymmetricalFirstStageLoad11 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=9e-6 W=197e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor12 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=9e-6 W=138e-6
mSecondStage1Transconductor13 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=9e-6 W=138e-6
mSymmetricalFirstStageLoad14 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=9e-6 W=197e-6
mMainBias15 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=15e-6
mSymmetricalFirstStageStageBias16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=317e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=70e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=34e-6
mSymmetricalFirstStageTransconductor19 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=64e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=322e-6
mSymmetricalFirstStageTransconductor21 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=64e-6
mMainBias22 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=52e-6
mMainBias23 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=27e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp149

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 1.20901 mW
** Area: 12957 (mu_m)^2
** Transit frequency: 3.38401 MHz
** Transit frequency with error factor: 3.38431 MHz
** Slew rate: 4.32116 V/mu_s
** Phase margin: 66.4632°
** CMRR: 152 dB
** negPSRR: 51 dB
** posPSRR: 67 dB
** VoutMax: 4.66001 V
** VoutMin: 0.330001 V
** VcmMax: 3.15001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.69211e+07 muA
** NormalTransistorPmos: -8.04699e+06 muA
** NormalTransistorPmos: -1.54749e+07 muA
** NormalTransistorNmos: 4.72411e+07 muA
** NormalTransistorNmos: 4.72401e+07 muA
** NormalTransistorNmos: 4.72411e+07 muA
** NormalTransistorNmos: 4.72401e+07 muA
** NormalTransistorPmos: -9.44839e+07 muA
** DiodeTransistorPmos: -9.44829e+07 muA
** NormalTransistorPmos: -4.72419e+07 muA
** NormalTransistorPmos: -4.72419e+07 muA
** NormalTransistorNmos: 4.34251e+07 muA
** NormalTransistorNmos: 4.34261e+07 muA
** NormalTransistorPmos: -4.34259e+07 muA
** NormalTransistorPmos: -4.34269e+07 muA
** DiodeTransistorPmos: -4.34259e+07 muA
** NormalTransistorNmos: 4.34251e+07 muA
** NormalTransistorNmos: 4.34261e+07 muA
** DiodeTransistorNmos: 8.04601e+06 muA
** DiodeTransistorNmos: 1.54741e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.69219e+07 muA


** Expected Voltages: 
** ibias: 3.35601  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 4.24901  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.737001  V
** outSourceVoltageBiasXXpXX1: 4.17901  V
** outVoltageBiasXXnXX0: 0.569001  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.172001  V
** innerTransistorStack2Load1: 0.172001  V
** sourceTransconductance: 3.26701  V
** innerStageBias: 4.40001  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V
** inner: 4.17601  V


.END