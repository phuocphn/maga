** Name: two_stage_single_output_op_amp_68_6

.MACRO two_stage_single_output_op_amp_68_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=130e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=9e-6 W=142e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=7e-6 W=142e-6
mMainBias5 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=3e-6 W=19e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=8e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=59e-6
mSecondStage1StageBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=397e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=81e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=145e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=145e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=334e-6
mSecondStage1Transconductor13 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=7e-6 W=221e-6
mFoldedCascodeFirstStageLoad14 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=81e-6
mMainBias15 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=14e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=9e-6 W=142e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=20e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=20e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=59e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mMainBias21 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
mSecondStage1StageBias22 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=3e-6 W=397e-6
mFoldedCascodeFirstStageLoad23 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=142e-6
mMainBias24 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=46e-6
mMainBias25 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=58e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_68_6

** Expected Performance Values: 
** Gain: 179 dB
** Power consumption: 1.80001 mW
** Area: 14951 (mu_m)^2
** Transit frequency: 2.69201 MHz
** Transit frequency with error factor: 2.69168 MHz
** Slew rate: 4.83295 V/mu_s
** Phase margin: 64.1713°
** CMRR: 136 dB
** VoutMax: 3.84001 V
** VoutMin: 0.430001 V
** VcmMax: 3.11001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.36201e+06 muA
** NormalTransistorPmos: -2.44309e+07 muA
** NormalTransistorPmos: -3.09899e+07 muA
** NormalTransistorNmos: 2.20401e+07 muA
** NormalTransistorNmos: 3.45221e+07 muA
** NormalTransistorNmos: 2.20401e+07 muA
** NormalTransistorNmos: 3.45221e+07 muA
** DiodeTransistorPmos: -2.20409e+07 muA
** NormalTransistorPmos: -2.20419e+07 muA
** NormalTransistorPmos: -2.20409e+07 muA
** DiodeTransistorPmos: -2.20419e+07 muA
** NormalTransistorPmos: -2.49669e+07 muA
** DiodeTransistorPmos: -2.49679e+07 muA
** NormalTransistorPmos: -1.24829e+07 muA
** NormalTransistorPmos: -1.24829e+07 muA
** NormalTransistorNmos: 2.12125e+08 muA
** NormalTransistorNmos: 2.12124e+08 muA
** NormalTransistorPmos: -2.12124e+08 muA
** DiodeTransistorPmos: -2.12123e+08 muA
** DiodeTransistorNmos: 2.44301e+07 muA
** DiodeTransistorNmos: 3.09891e+07 muA
** DiodeTransistorPmos: -3.36299e+06 muA
** NormalTransistorPmos: -3.36399e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.27401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.43601  V
** outSourceVoltageBiasXXpXX1: 4.21801  V
** outSourceVoltageBiasXXpXX2: 4.13801  V
** outVoltageBiasXXnXX1: 0.905001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.15501  V
** innerTransistorStack2Load2: 4.15601  V
** out1: 3.34501  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.38701  V
** innerTransconductance: 0.217001  V
** inner: 4.21601  V
** inner: 4.13401  V


.END