** Name: two_stage_single_output_op_amp_1_5

.MACRO two_stage_single_output_op_amp_1_5 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=150e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=13e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=48e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=163e-6
mSimpleFirstStageLoad7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=150e-6
mMainBias8 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=44e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=43e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=97e-6
mMainBias11 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=13e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=48e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=43e-6
mMainBias14 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_1_5

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 1.53601 mW
** Area: 4035 (mu_m)^2
** Transit frequency: 4.12701 MHz
** Transit frequency with error factor: 4.10375 MHz
** Slew rate: 6.35057 V/mu_s
** Phase margin: 65.3172°
** CMRR: 88 dB
** negPSRR: 90 dB
** posPSRR: 200 dB
** VoutMax: 3.23001 V
** VoutMin: 0.150001 V
** VcmMax: 3.44001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 4.25181e+07 muA
** NormalTransistorPmos: -6.75999e+06 muA
** DiodeTransistorNmos: 4.09861e+07 muA
** NormalTransistorNmos: 4.09861e+07 muA
** NormalTransistorPmos: -8.19729e+07 muA
** NormalTransistorPmos: -4.09869e+07 muA
** NormalTransistorPmos: -4.09869e+07 muA
** NormalTransistorNmos: 1.55887e+08 muA
** NormalTransistorPmos: -1.55886e+08 muA
** DiodeTransistorPmos: -1.55887e+08 muA
** DiodeTransistorNmos: 6.75901e+06 muA
** DiodeTransistorPmos: -4.25189e+07 muA
** NormalTransistorPmos: -4.25199e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.66201  V
** outSourceVoltageBiasXXpXX1: 3.83101  V
** outVoltageBiasXXnXX0: 0.687001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceTransconductance: 3.75401  V
** inner: 3.82801  V


.END