** Name: two_stage_single_output_op_amp_123_8

.MACRO two_stage_single_output_op_amp_123_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=7e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=20e-6
mMainBias3 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mTelescopicFirstStageLoad4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=10e-6 W=145e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=10e-6 W=145e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=50e-6
mTelescopicFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=116e-6
mTelescopicFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=20e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=10e-6 W=67e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=10e-6 W=67e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=158e-6
mTelescopicFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=20e-6
mMainBias14 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=30e-6
mTelescopicFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=10e-6 W=145e-6
mMainBias17 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=492e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=406e-6
mTelescopicFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=10e-6 W=145e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.6001e-12
.EOM two_stage_single_output_op_amp_123_8

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 2.46201 mW
** Area: 14998 (mu_m)^2
** Transit frequency: 2.54201 MHz
** Transit frequency with error factor: 2.54223 MHz
** Slew rate: 7.20989 V/mu_s
** Phase margin: 60.1606°
** CMRR: 142 dB
** VoutMax: 4.53001 V
** VoutMin: 0.860001 V
** VcmMax: 3.68001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorNmos: 5.23201e+06 muA
** NormalTransistorPmos: -5.12789e+07 muA
** NormalTransistorNmos: 1.27601e+07 muA
** NormalTransistorNmos: 1.27601e+07 muA
** DiodeTransistorPmos: -1.27609e+07 muA
** NormalTransistorPmos: -1.27619e+07 muA
** NormalTransistorPmos: -1.27609e+07 muA
** DiodeTransistorPmos: -1.27619e+07 muA
** NormalTransistorNmos: 7.67991e+07 muA
** NormalTransistorNmos: 7.67981e+07 muA
** NormalTransistorNmos: 1.27611e+07 muA
** NormalTransistorNmos: 1.27611e+07 muA
** NormalTransistorNmos: 4.00319e+08 muA
** NormalTransistorNmos: 4.00318e+08 muA
** NormalTransistorPmos: -4.00318e+08 muA
** DiodeTransistorNmos: 5.12781e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.23299e+06 muA


** Expected Voltages: 
** ibias: 1.18701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.65001  V
** out: 2.5  V
** outFirstStage: 3.96401  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX0: 4.24801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.21301  V
** innerStageBias: 0.482001  V
** innerTransistorStack1Load2: 4.21101  V
** out1: 3.42601  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.482001  V


.END