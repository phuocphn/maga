** Name: two_stage_single_output_op_amp_206_7

.MACRO two_stage_single_output_op_amp_206_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=9e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=82e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=37e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=31e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=20e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=8e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=45e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=37e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=82e-6
mSecondStage1StageBias12 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=258e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=9e-6 W=10e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=45e-6
mSimpleFirstStageLoad15 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=229e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=36e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=36e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=257e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=229e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=30e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=125e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_206_7

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 8.04901 mW
** Area: 7435 (mu_m)^2
** Transit frequency: 3.96301 MHz
** Transit frequency with error factor: 3.96134 MHz
** Slew rate: 3.73455 V/mu_s
** Phase margin: 65.3172°
** CMRR: 110 dB
** VoutMax: 4.25 V
** VoutMin: 0.690001 V
** VcmMax: 4.76001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorPmos: -3.81789e+07 muA
** NormalTransistorPmos: -1.56834e+08 muA
** DiodeTransistorNmos: 3.64921e+07 muA
** NormalTransistorNmos: 3.64931e+07 muA
** NormalTransistorNmos: 3.64941e+07 muA
** DiodeTransistorNmos: 3.64931e+07 muA
** NormalTransistorPmos: -4.50639e+07 muA
** NormalTransistorPmos: -4.50649e+07 muA
** NormalTransistorPmos: -4.50659e+07 muA
** NormalTransistorPmos: -4.50649e+07 muA
** NormalTransistorNmos: 1.71411e+07 muA
** DiodeTransistorNmos: 1.71401e+07 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 1.30472e+09 muA
** NormalTransistorPmos: -1.30471e+09 muA
** DiodeTransistorNmos: 3.81781e+07 muA
** NormalTransistorNmos: 3.81771e+07 muA
** DiodeTransistorNmos: 1.56835e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.12201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.14001  V
** outSourceVoltageBiasXXnXX1: 0.570001  V
** outSourceVoltageBiasXXpXX1: 3.97601  V
** outVoltageBiasXXnXX2: 1.09301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.06401  V
** innerTransistorStack1Load1: 1.06501  V
** innerTransistorStack1Load2: 3.86701  V
** innerTransistorStack2Load2: 3.86701  V
** sourceTransconductance: 1.94501  V
** inner: 0.569001  V


.END