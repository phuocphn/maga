** Name: two_stage_single_output_op_amp_34_11

.MACRO two_stage_single_output_op_amp_34_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=498e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=25e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=193e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=51e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=60e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=25e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=556e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=498e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=140e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=60e-6
mMainBias14 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=23e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=104e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=193e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=522e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=5e-6 W=600e-6
mSimpleFirstStageLoad19 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=5e-6 W=111e-6
mMainBias20 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=370e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.10001e-12
.EOM two_stage_single_output_op_amp_34_11

** Expected Performance Values: 
** Gain: 144 dB
** Power consumption: 6.82101 mW
** Area: 14777 (mu_m)^2
** Transit frequency: 4.84601 MHz
** Transit frequency with error factor: 4.84408 MHz
** Slew rate: 4.5669 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** negPSRR: 103 dB
** posPSRR: 98 dB
** VoutMax: 4.25 V
** VoutMin: 0.860001 V
** VcmMax: 4.47001 V
** VcmMin: 1.51001 V


** Expected Currents: 
** NormalTransistorNmos: 2.28411e+07 muA
** NormalTransistorNmos: 1.03564e+08 muA
** NormalTransistorPmos: -6.40508e+08 muA
** DiodeTransistorPmos: -1.63269e+07 muA
** NormalTransistorPmos: -1.63269e+07 muA
** NormalTransistorPmos: -1.63269e+07 muA
** NormalTransistorNmos: 3.26511e+07 muA
** DiodeTransistorNmos: 3.26501e+07 muA
** NormalTransistorNmos: 1.63261e+07 muA
** NormalTransistorNmos: 1.63261e+07 muA
** NormalTransistorNmos: 5.54589e+08 muA
** NormalTransistorNmos: 5.54588e+08 muA
** NormalTransistorPmos: -5.54588e+08 muA
** NormalTransistorPmos: -5.54589e+08 muA
** DiodeTransistorNmos: 6.40509e+08 muA
** NormalTransistorNmos: 6.40509e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.28419e+07 muA
** DiodeTransistorPmos: -1.03563e+08 muA


** Expected Voltages: 
** ibias: 1.18001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.19201  V
** outInputVoltageBiasXXnXX1: 1.36401  V
** outSourceVoltageBiasXXnXX1: 0.682001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX0: 4.12401  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.45201  V
** out1: 4.26701  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.468001  V
** innerTransconductance: 4.75601  V
** inner: 0.682001  V


.END