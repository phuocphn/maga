** Name: two_stage_single_output_op_amp_129_1

.MACRO two_stage_single_output_op_amp_129_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=178e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=10e-6 W=62e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSimpleFirstStageLoad4 FirstStageYout1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=72e-6
mSecondStage1Transconductor5 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=415e-6
mSimpleFirstStageLoad6 outFirstStage inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=72e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=183e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=10e-6 W=62e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=174e-6
mMainBias10 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=564e-6
mSecondStage1StageBias11 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=31e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=183e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.4001e-12
.EOM two_stage_single_output_op_amp_129_1

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 3.64801 mW
** Area: 8685 (mu_m)^2
** Transit frequency: 3.39601 MHz
** Transit frequency with error factor: 3.38851 MHz
** Slew rate: 4.58532 V/mu_s
** Phase margin: 60.1606°
** CMRR: 84 dB
** VoutMax: 4.84001 V
** VoutMin: 0.150001 V
** VcmMax: 4.07001 V
** VcmMin: -0.159999 V


** Expected Currents: 
** NormalTransistorPmos: -2.44701e+08 muA
** NormalTransistorPmos: -6.29509e+07 muA
** NormalTransistorPmos: -6.29509e+07 muA
** DiodeTransistorPmos: -6.29509e+07 muA
** NormalTransistorNmos: 1.00702e+08 muA
** NormalTransistorNmos: 1.00702e+08 muA
** NormalTransistorPmos: -7.55029e+07 muA
** NormalTransistorPmos: -3.77509e+07 muA
** NormalTransistorPmos: -3.77509e+07 muA
** NormalTransistorNmos: 2.63568e+08 muA
** NormalTransistorPmos: -2.63565e+08 muA
** DiodeTransistorNmos: 2.44702e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.810001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.68601  V
** out1: 2.37201  V
** sourceTransconductance: 3.27801  V


.END