** Name: two_stage_single_output_op_amp_108_9

.MACRO two_stage_single_output_op_amp_108_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=28e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=13e-6
mTelescopicFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=518e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=147e-6
mTelescopicFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=138e-6
mTelescopicFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=138e-6
mTelescopicFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=86e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=86e-6
mMainBias14 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=123e-6
mTelescopicFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=46e-6
mTelescopicFirstStageTransconductor16 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=176e-6
mTelescopicFirstStageTransconductor17 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=176e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=13e-6
mMainBias19 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=25e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=10e-6 W=361e-6
mTelescopicFirstStageLoad21 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=46e-6
mMainBias22 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=18e-6
mMainBias23 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=56e-6
mTelescopicFirstStageStageBias24 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=518e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.3001e-12
.EOM two_stage_single_output_op_amp_108_9

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 14.0451 mW
** Area: 14997 (mu_m)^2
** Transit frequency: 2.91101 MHz
** Transit frequency with error factor: 2.91083 MHz
** Slew rate: 30.3088 V/mu_s
** Phase margin: 60.1606°
** CMRR: 129 dB
** VoutMax: 3.10001 V
** VoutMin: 1 V
** VcmMax: 3.01001 V
** VcmMin: -0.0699999 V


** Expected Currents: 
** NormalTransistorNmos: 3.37927e+08 muA
** NormalTransistorPmos: -1.40099e+07 muA
** NormalTransistorPmos: -1.91169e+07 muA
** NormalTransistorPmos: -4.30949e+07 muA
** NormalTransistorPmos: -3.30839e+07 muA
** NormalTransistorPmos: -3.30839e+07 muA
** NormalTransistorNmos: 3.30831e+07 muA
** NormalTransistorNmos: 3.30821e+07 muA
** NormalTransistorNmos: 3.30831e+07 muA
** NormalTransistorNmos: 3.30821e+07 muA
** NormalTransistorPmos: -4.04095e+08 muA
** DiodeTransistorPmos: -4.04094e+08 muA
** NormalTransistorPmos: -3.30849e+07 muA
** NormalTransistorPmos: -3.30849e+07 muA
** NormalTransistorNmos: 2.30864e+09 muA
** DiodeTransistorNmos: 2.30864e+09 muA
** NormalTransistorPmos: -2.30863e+09 muA
** DiodeTransistorNmos: 1.40091e+07 muA
** DiodeTransistorNmos: 1.91161e+07 muA
** NormalTransistorNmos: 1.91151e+07 muA
** DiodeTransistorNmos: 4.30941e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -3.37926e+08 muA


** Expected Voltages: 
** ibias: 3.28201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.41001  V
** out: 2.5  V
** outFirstStage: 2.53501  V
** outSourceVoltageBiasXXnXX1: 0.705001  V
** outSourceVoltageBiasXXpXX1: 4.14201  V
** outVoltageBiasXXnXX0: 0.661001  V
** outVoltageBiasXXnXX2: 0.705001  V
** outVoltageBiasXXpXX2: 2.14601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.33401  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.05601  V
** sourceGCC2: 3.05601  V
** inner: 0.705001  V
** inner: 4.13801  V


.END