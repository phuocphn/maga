** Name: two_stage_single_output_op_amp_82_9

.MACRO two_stage_single_output_op_amp_82_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=29e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=184e-6
mMainBias4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=9e-6 W=26e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=63e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=215e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=7e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=7e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=63e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=184e-6
mMainBias14 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=26e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=9e-6 W=215e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=29e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=162e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=105e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=105e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=336e-6
mFoldedCascodeFirstStageLoad21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=162e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=239e-6
mMainBias23 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=104e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_82_9

** Expected Performance Values: 
** Gain: 117 dB
** Power consumption: 7.13701 mW
** Area: 7856 (mu_m)^2
** Transit frequency: 4.98601 MHz
** Transit frequency with error factor: 4.98587 MHz
** Slew rate: 13.2789 V/mu_s
** Phase margin: 60.1606°
** CMRR: 137 dB
** VoutMax: 4.25 V
** VoutMin: 1.70001 V
** VcmMax: 5.17001 V
** VcmMin: 1.68001 V


** Expected Currents: 
** NormalTransistorPmos: -2.38166e+08 muA
** NormalTransistorPmos: -1.03403e+08 muA
** NormalTransistorPmos: -6.57939e+07 muA
** NormalTransistorPmos: -1.06456e+08 muA
** NormalTransistorPmos: -6.57939e+07 muA
** NormalTransistorPmos: -1.06456e+08 muA
** DiodeTransistorNmos: 6.57931e+07 muA
** NormalTransistorNmos: 6.57921e+07 muA
** NormalTransistorNmos: 6.57931e+07 muA
** DiodeTransistorNmos: 6.57921e+07 muA
** NormalTransistorNmos: 8.13231e+07 muA
** DiodeTransistorNmos: 8.13221e+07 muA
** NormalTransistorNmos: 4.06621e+07 muA
** NormalTransistorNmos: 4.06621e+07 muA
** NormalTransistorNmos: 8.52886e+08 muA
** DiodeTransistorNmos: 8.52885e+08 muA
** NormalTransistorPmos: -8.52885e+08 muA
** DiodeTransistorNmos: 2.38167e+08 muA
** NormalTransistorNmos: 2.38166e+08 muA
** DiodeTransistorNmos: 1.03404e+08 muA
** NormalTransistorNmos: 1.03403e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.15801  V
** outInputVoltageBiasXXnXX2: 2.10401  V
** outSourceVoltageBiasXXnXX1: 0.579001  V
** outSourceVoltageBiasXXnXX2: 1.05201  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.687001  V
** innerTransistorStack2Load2: 0.688001  V
** out1: 1.25601  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.56901  V
** inner: 0.578001  V
** inner: 1.04601  V


.END