** Name: symmetrical_op_amp51

.MACRO symmetrical_op_amp51 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=28e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=27e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=25e-6
mSymmetricalFirstStageLoad4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=27e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=24e-6
mMainBias6 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=32e-6
mSymmetricalFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=93e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=79e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=79e-6
mMainBias10 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=264e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=5e-6 W=33e-6
mSecondStage1Transconductor12 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=33e-6
mSymmetricalFirstStageStageBias13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=93e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=240e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias15 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=240e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=24e-6
mMainBias17 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=354e-6
mSymmetricalFirstStageTransconductor18 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=69e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias19 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=3e-6 W=45e-6
mMainBias20 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=24e-6
mSecondStage1StageBias21 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=94e-6
mSymmetricalFirstStageTransconductor22 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=69e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp51

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 2.19401 mW
** Area: 8016 (mu_m)^2
** Transit frequency: 2.95501 MHz
** Transit frequency with error factor: 2.95509 MHz
** Slew rate: 5.67008 V/mu_s
** Phase margin: 68.182°
** CMRR: 138 dB
** negPSRR: 46 dB
** posPSRR: 57 dB
** VoutMax: 4.48001 V
** VoutMin: 0.560001 V
** VcmMax: 3.03001 V
** VcmMin: 0.0900001 V


** Expected Currents: 
** NormalTransistorNmos: 1.0707e+08 muA
** NormalTransistorPmos: -1.01399e+07 muA
** NormalTransistorPmos: -1.48769e+08 muA
** DiodeTransistorNmos: 1.96471e+07 muA
** DiodeTransistorNmos: 1.96471e+07 muA
** NormalTransistorPmos: -3.92959e+07 muA
** DiodeTransistorPmos: -3.92949e+07 muA
** NormalTransistorPmos: -1.96479e+07 muA
** NormalTransistorPmos: -1.96479e+07 muA
** NormalTransistorNmos: 5.67761e+07 muA
** NormalTransistorNmos: 5.67771e+07 muA
** NormalTransistorPmos: -5.67769e+07 muA
** NormalTransistorPmos: -5.67779e+07 muA
** NormalTransistorPmos: -5.67769e+07 muA
** NormalTransistorPmos: -5.67779e+07 muA
** NormalTransistorNmos: 5.67761e+07 muA
** NormalTransistorNmos: 5.67771e+07 muA
** DiodeTransistorNmos: 1.01391e+07 muA
** DiodeTransistorNmos: 1.4877e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.07069e+08 muA


** Expected Voltages: 
** ibias: 3.34001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 3.68601  V
** inOutputTransconductanceComplementarySecondStage: 0.968001  V
** inSourceTransconductanceComplementarySecondStage: 0.650001  V
** innerComplementarySecondStage: 4.23601  V
** inputVoltageBiasXXnXX0: 0.559001  V
** out: 2.5  V
** outFirstStage: 0.650001  V
** outSourceVoltageBiasXXpXX1: 4.17101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.37201  V
** innerStageBias: 4.56701  V
** innerTransconductance: 0.245001  V
** inner: 4.70801  V
** inner: 0.245001  V
** inner: 4.16801  V


.END