** Name: one_stage_single_output_op_amp78

.MACRO one_stage_single_output_op_amp78 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=74e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
mMainBias3 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=45e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=9e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=84e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=79e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=79e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=45e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias12 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mFoldedCascodeFirstStageLoad13 out FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=74e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerOutputLoad2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=351e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=291e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=291e-6
mFoldedCascodeFirstStageLoad17 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=351e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp78

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 1.29201 mW
** Area: 4554 (mu_m)^2
** Transit frequency: 2.97601 MHz
** Transit frequency with error factor: 2.97553 MHz
** Slew rate: 3.5455 V/mu_s
** Phase margin: 86.5167°
** CMRR: 147 dB
** VoutMax: 4.08001 V
** VoutMin: 0.760001 V
** VcmMax: 5.20001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 3.18451e+07 muA
** NormalTransistorPmos: -7.12739e+07 muA
** NormalTransistorPmos: -1.08238e+08 muA
** NormalTransistorPmos: -7.12759e+07 muA
** NormalTransistorPmos: -1.0824e+08 muA
** DiodeTransistorNmos: 7.12731e+07 muA
** DiodeTransistorNmos: 7.12741e+07 muA
** NormalTransistorNmos: 7.12751e+07 muA
** NormalTransistorNmos: 7.12741e+07 muA
** NormalTransistorNmos: 7.39291e+07 muA
** DiodeTransistorNmos: 7.39301e+07 muA
** NormalTransistorNmos: 3.69641e+07 muA
** NormalTransistorNmos: 3.69641e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.18459e+07 muA
** DiodeTransistorPmos: -3.18469e+07 muA


** Expected Voltages: 
** ibias: 1.20501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.603001  V
** outSourceVoltageBiasXXpXX1: 4.23101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.16801  V
** innerTransistorStack1Load2: 0.612001  V
** innerTransistorStack2Load2: 0.612001  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.89801  V
** inner: 0.601001  V


.END