** Name: two_stage_single_output_op_amp_144_9

.MACRO two_stage_single_output_op_amp_144_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=11e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=137e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=23e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=11e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=137e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=76e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=600e-6
mMainBias17 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=59e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=216e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=600e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=36e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_144_9

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 10.3131 mW
** Area: 5222 (mu_m)^2
** Transit frequency: 3.42301 MHz
** Transit frequency with error factor: 3.41939 MHz
** Slew rate: 3.6639 V/mu_s
** Phase margin: 66.4632°
** CMRR: 126 dB
** VoutMax: 4.25 V
** VoutMin: 1.40001 V
** VcmMax: 4.93001 V
** VcmMin: 1 V


** Expected Currents: 
** NormalTransistorPmos: -5.87859e+07 muA
** NormalTransistorPmos: -3.60259e+07 muA
** NormalTransistorNmos: 5.99728e+08 muA
** NormalTransistorNmos: 5.99727e+08 muA
** DiodeTransistorNmos: 5.99728e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** NormalTransistorPmos: -6.08325e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** NormalTransistorNmos: 1.71971e+07 muA
** NormalTransistorNmos: 8.59901e+06 muA
** NormalTransistorNmos: 8.59901e+06 muA
** NormalTransistorNmos: 7.31045e+08 muA
** DiodeTransistorNmos: 7.31044e+08 muA
** NormalTransistorPmos: -7.31044e+08 muA
** DiodeTransistorNmos: 5.87851e+07 muA
** NormalTransistorNmos: 5.87841e+07 muA
** DiodeTransistorNmos: 3.60251e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.81001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.905001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.833001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.940001  V
** innerTransistorStack1Load2: 4.21001  V
** innerTransistorStack2Load2: 4.21001  V
** out1: 2.09501  V
** sourceTransconductance: 1.92401  V
** inner: 0.900001  V


.END