** Name: two_stage_single_output_op_amp_59_2

.MACRO two_stage_single_output_op_amp_59_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=144e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=103e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=18e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=97e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=408e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=408e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=276e-6
mMainBias10 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=574e-6
mSecondStage1Transconductor11 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=406e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=97e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=194e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=103e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=62e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=62e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=266e-6
mMainBias18 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=66e-6
mSecondStage1StageBias19 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=466e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=4e-6 W=104e-6
mMainBias21 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=83e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.2001e-12
.EOM two_stage_single_output_op_amp_59_2

** Expected Performance Values: 
** Gain: 135 dB
** Power consumption: 4.03901 mW
** Area: 14997 (mu_m)^2
** Transit frequency: 3.85901 MHz
** Transit frequency with error factor: 3.85902 MHz
** Slew rate: 5.29759 V/mu_s
** Phase margin: 60.1606°
** CMRR: 129 dB
** VoutMax: 4.75 V
** VoutMin: 0.300001 V
** VcmMax: 3.16001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.82761e+08 muA
** NormalTransistorPmos: -3.72289e+07 muA
** NormalTransistorPmos: -4.58919e+07 muA
** NormalTransistorNmos: 7.55511e+07 muA
** NormalTransistorNmos: 1.29516e+08 muA
** NormalTransistorNmos: 7.55501e+07 muA
** NormalTransistorNmos: 1.29516e+08 muA
** NormalTransistorPmos: -7.55519e+07 muA
** NormalTransistorPmos: -7.55509e+07 muA
** DiodeTransistorPmos: -7.55519e+07 muA
** NormalTransistorPmos: -1.07928e+08 muA
** NormalTransistorPmos: -1.07929e+08 muA
** NormalTransistorPmos: -5.39639e+07 muA
** NormalTransistorPmos: -5.39639e+07 muA
** NormalTransistorNmos: 2.62839e+08 muA
** NormalTransistorNmos: 2.6284e+08 muA
** NormalTransistorPmos: -2.62838e+08 muA
** DiodeTransistorNmos: 3.72281e+07 muA
** DiodeTransistorNmos: 4.58911e+07 muA
** DiodeTransistorPmos: -1.8276e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.921001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.02901  V
** innerStageBias: 4.40001  V
** out1: 3.06001  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.375  V
** innerTransconductance: 0.364001  V


.END