** Name: two_stage_single_output_op_amp_116_9

.MACRO two_stage_single_output_op_amp_116_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=7e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=12e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=499e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=210e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=36e-6
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=141e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=15e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=29e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=29e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=29e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=12e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mMainBias13 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSecondStage1StageBias14 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=210e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=29e-6
mTelescopicFirstStageStageBias16 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=499e-6
mTelescopicFirstStageLoad17 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=141e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=161e-6
mTelescopicFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=32e-6
mMainBias20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=6e-6
mMainBias21 outVoltageBiasXXnXX3 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=179e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.7001e-12
.EOM two_stage_single_output_op_amp_116_9

** Expected Performance Values: 
** Gain: 148 dB
** Power consumption: 2.04301 mW
** Area: 14983 (mu_m)^2
** Transit frequency: 2.50101 MHz
** Transit frequency with error factor: 2.50076 MHz
** Slew rate: 8.1505 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.68001 V
** VoutMin: 0.920001 V
** VcmMax: 4.37001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 5.73501e+06 muA
** NormalTransistorPmos: -2.28699e+06 muA
** NormalTransistorPmos: -6.78889e+07 muA
** NormalTransistorNmos: 1.38091e+07 muA
** NormalTransistorNmos: 1.38091e+07 muA
** NormalTransistorPmos: -1.38099e+07 muA
** NormalTransistorPmos: -1.38099e+07 muA
** DiodeTransistorPmos: -1.38099e+07 muA
** NormalTransistorNmos: 9.55051e+07 muA
** DiodeTransistorNmos: 9.55041e+07 muA
** NormalTransistorNmos: 1.38091e+07 muA
** NormalTransistorNmos: 1.38091e+07 muA
** NormalTransistorNmos: 2.95165e+08 muA
** DiodeTransistorNmos: 2.95166e+08 muA
** NormalTransistorPmos: -2.95164e+08 muA
** DiodeTransistorNmos: 2.28601e+06 muA
** NormalTransistorNmos: 2.28601e+06 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 6.78881e+07 muA
** DiodeTransistorPmos: -5.73599e+06 muA


** Expected Voltages: 
** ibias: 1.32601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.14401  V
** out: 2.5  V
** outFirstStage: 4.11501  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.664001  V
** outVoltageBiasXXnXX3: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.27001  V
** out1: 3.55101  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.555001  V
** inner: 0.660001  V


.END