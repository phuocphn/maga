** Name: two_stage_single_output_op_amp_78_7

.MACRO two_stage_single_output_op_amp_78_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=66e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=8e-6 W=35e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=150e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=16e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=45e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=8e-6 W=35e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=17e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=16e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=150e-6
mSecondStage1StageBias13 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=224e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=66e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerOutputLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=206e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=39e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=159e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=213e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_78_7

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 7.43901 mW
** Area: 7159 (mu_m)^2
** Transit frequency: 3.88801 MHz
** Transit frequency with error factor: 3.8884 MHz
** Slew rate: 3.50036 V/mu_s
** Phase margin: 71.0468°
** CMRR: 149 dB
** VoutMax: 4.25 V
** VoutMin: 0.670001 V
** VcmMax: 5.17001 V
** VcmMin: 1.55001 V


** Expected Currents: 
** NormalTransistorPmos: -1.59452e+08 muA
** NormalTransistorPmos: -2.13976e+08 muA
** NormalTransistorPmos: -1.58389e+07 muA
** NormalTransistorPmos: -2.43329e+07 muA
** NormalTransistorPmos: -1.58389e+07 muA
** NormalTransistorPmos: -2.43329e+07 muA
** DiodeTransistorNmos: 1.58381e+07 muA
** DiodeTransistorNmos: 1.58371e+07 muA
** NormalTransistorNmos: 1.58381e+07 muA
** NormalTransistorNmos: 1.58371e+07 muA
** NormalTransistorNmos: 1.69851e+07 muA
** DiodeTransistorNmos: 1.69841e+07 muA
** NormalTransistorNmos: 8.49301e+06 muA
** NormalTransistorNmos: 8.49301e+06 muA
** NormalTransistorNmos: 1.04581e+09 muA
** NormalTransistorPmos: -1.0458e+09 muA
** DiodeTransistorNmos: 1.59453e+08 muA
** NormalTransistorNmos: 1.59452e+08 muA
** DiodeTransistorNmos: 2.13977e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.40001  V
** outSourceVoltageBiasXXnXX1: 0.700001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 1.07201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.16601  V
** innerTransistorStack1Load2: 0.611001  V
** innerTransistorStack2Load2: 0.610001  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.94101  V
** inner: 0.698001  V


.END