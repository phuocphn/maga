** Name: two_stage_single_output_op_amp_189_9

.MACRO two_stage_single_output_op_amp_189_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=42e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=4e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=17e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=414e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=75e-6
mSimpleFirstStageLoad10 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=42e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=31e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=17e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=414e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=1e-6 W=14e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=75e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=349e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=349e-6
mSimpleFirstStageLoad18 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=596e-6
mMainBias19 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=269e-6
mSimpleFirstStageLoad21 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=596e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=55e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_189_9

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 10.8561 mW
** Area: 5405 (mu_m)^2
** Transit frequency: 7.16601 MHz
** Transit frequency with error factor: 7.16138 MHz
** Slew rate: 6.75375 V/mu_s
** Phase margin: 64.7443°
** CMRR: 124 dB
** VoutMax: 4.25 V
** VoutMin: 0.800001 V
** VcmMax: 4.99001 V
** VcmMin: 1.55001 V


** Expected Currents: 
** NormalTransistorPmos: -5.53649e+07 muA
** NormalTransistorPmos: -2.68329e+07 muA
** NormalTransistorNmos: 3.35847e+08 muA
** NormalTransistorNmos: 3.35848e+08 muA
** DiodeTransistorNmos: 3.35847e+08 muA
** NormalTransistorPmos: -3.51718e+08 muA
** NormalTransistorPmos: -3.51719e+08 muA
** NormalTransistorPmos: -3.51719e+08 muA
** NormalTransistorPmos: -3.51719e+08 muA
** NormalTransistorNmos: 3.17431e+07 muA
** NormalTransistorNmos: 3.17421e+07 muA
** NormalTransistorNmos: 1.58721e+07 muA
** NormalTransistorNmos: 1.58721e+07 muA
** NormalTransistorNmos: 1.36564e+09 muA
** DiodeTransistorNmos: 1.36564e+09 muA
** NormalTransistorPmos: -1.36563e+09 muA
** DiodeTransistorNmos: 5.53641e+07 muA
** NormalTransistorNmos: 5.53631e+07 muA
** DiodeTransistorNmos: 2.68321e+07 muA
** DiodeTransistorNmos: 2.68311e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.69501  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.20401  V
** outSourceVoltageBiasXXnXX1: 0.602001  V
** outSourceVoltageBiasXXnXX2: 0.804001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 1.09901  V
** innerTransistorStack1Load2: 4.15401  V
** innerTransistorStack2Load2: 4.15401  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 0.602001  V


.END