** Name: symmetrical_op_amp8

.MACRO symmetrical_op_amp8 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=9e-6 W=54e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=5e-6 W=36e-6
mSecondStage1Transconductor10 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=36e-6
mSymmetricalFirstStageStageBias11 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=9e-6 W=129e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mMainBias13 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=9e-6 W=89e-6
mSymmetricalFirstStageTransconductor14 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=62e-6
mSecondStage1StageBias15 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=89e-6
mSymmetricalFirstStageTransconductor16 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=62e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp8

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 0.664001 mW
** Area: 3582 (mu_m)^2
** Transit frequency: 2.76101 MHz
** Transit frequency with error factor: 2.76149 MHz
** Slew rate: 3.58566 V/mu_s
** Phase margin: 85.3708°
** CMRR: 148 dB
** negPSRR: 50 dB
** posPSRR: 64 dB
** VoutMax: 3.98001 V
** VoutMin: 0.440001 V
** VcmMax: 3.92001 V
** VcmMin: 0.0400001 V


** Expected Currents: 
** NormalTransistorPmos: -1.67129e+07 muA
** DiodeTransistorNmos: 1.21111e+07 muA
** DiodeTransistorNmos: 1.21111e+07 muA
** NormalTransistorPmos: -2.42249e+07 muA
** NormalTransistorPmos: -1.21119e+07 muA
** NormalTransistorPmos: -1.21119e+07 muA
** NormalTransistorNmos: 3.59081e+07 muA
** NormalTransistorNmos: 3.59091e+07 muA
** NormalTransistorPmos: -3.59089e+07 muA
** NormalTransistorPmos: -3.59099e+07 muA
** DiodeTransistorPmos: -3.59109e+07 muA
** DiodeTransistorPmos: -3.59119e+07 muA
** NormalTransistorNmos: 3.59101e+07 muA
** NormalTransistorNmos: 3.59091e+07 muA
** DiodeTransistorNmos: 1.67121e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.849001  V
** inSourceStageBiasComplementarySecondStage: 4.12601  V
** inSourceTransconductanceComplementarySecondStage: 0.607001  V
** innerComplementarySecondStage: 3.11201  V
** out: 2.5  V
** outFirstStage: 0.607001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.27301  V
** innerStageBias: 3.82601  V
** innerTransconductance: 0.202001  V
** inner: 0.202001  V


.END