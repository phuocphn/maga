** Name: two_stage_single_output_op_amp_23_1

.MACRO two_stage_single_output_op_amp_23_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=6e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=137e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=244e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=81e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=81e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=81e-6
mMainBias8 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=187e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=504e-6
mSimpleFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=81e-6
mSimpleFirstStageTransconductor11 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=66e-6
mSimpleFirstStageStageBias12 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=145e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=6e-6 W=161e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mSecondStage1StageBias15 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=66e-6
mMainBias17 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=515e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_23_1

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 5.30501 mW
** Area: 7019 (mu_m)^2
** Transit frequency: 7.34901 MHz
** Transit frequency with error factor: 7.34263 MHz
** Slew rate: 8.35549 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** negPSRR: 106 dB
** posPSRR: 221 dB
** VoutMax: 4.83001 V
** VoutMin: 0.150001 V
** VcmMax: 3.12001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.62106e+08 muA
** NormalTransistorPmos: -2.69652e+08 muA
** NormalTransistorPmos: -1.15439e+07 muA
** NormalTransistorNmos: 3.86231e+07 muA
** NormalTransistorNmos: 3.86221e+07 muA
** NormalTransistorNmos: 3.86211e+07 muA
** NormalTransistorNmos: 3.86221e+07 muA
** NormalTransistorPmos: -7.72429e+07 muA
** NormalTransistorPmos: -7.72439e+07 muA
** NormalTransistorPmos: -3.86219e+07 muA
** NormalTransistorPmos: -3.86219e+07 muA
** NormalTransistorNmos: 3.20403e+08 muA
** NormalTransistorPmos: -3.20402e+08 muA
** DiodeTransistorNmos: 2.69653e+08 muA
** DiodeTransistorNmos: 1.15431e+07 muA
** DiodeTransistorPmos: -3.62105e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXpXX1: 3.72701  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.557001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerStageBias: 4.69101  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.24501  V


.END