** Name: two_stage_single_output_op_amp_159_1

.MACRO two_stage_single_output_op_amp_159_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=15e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
mMainBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mSimpleFirstStageLoad5 FirstStageYout1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=170e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=586e-6
mSimpleFirstStageLoad7 outFirstStage ibias sourceNmos sourceNmos nmos4 L=5e-6 W=170e-6
mMainBias8 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=111e-6
mMainBias9 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=68e-6
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=104e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=530e-6
mSimpleFirstStageLoad12 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=304e-6
mSecondStage1StageBias14 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=558e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=15e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=530e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.5e-12
.EOM two_stage_single_output_op_amp_159_1

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 7.34201 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 4.84401 MHz
** Transit frequency with error factor: 4.84047 MHz
** Slew rate: 10.1055 V/mu_s
** Phase margin: 60.1606°
** CMRR: 70 dB
** VoutMax: 4.66001 V
** VoutMin: 0.150001 V
** VcmMax: 3.01001 V
** VcmMin: -0.369999 V


** Expected Currents: 
** NormalTransistorNmos: 7.39701e+07 muA
** NormalTransistorNmos: 4.48311e+07 muA
** NormalTransistorPmos: -7.31399e+06 muA
** NormalTransistorPmos: -7.31399e+06 muA
** DiodeTransistorPmos: -7.31399e+06 muA
** NormalTransistorNmos: 1.11717e+08 muA
** NormalTransistorNmos: 1.11717e+08 muA
** NormalTransistorPmos: -2.08806e+08 muA
** NormalTransistorPmos: -2.08807e+08 muA
** NormalTransistorPmos: -1.04402e+08 muA
** NormalTransistorPmos: -1.04402e+08 muA
** NormalTransistorNmos: 1.11612e+09 muA
** NormalTransistorPmos: -1.11611e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.39709e+07 muA
** DiodeTransistorPmos: -4.48319e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXpXX1: 3.84601  V
** outVoltageBiasXXpXX2: 4.10001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.79401  V
** innerStageBias: 4.60601  V
** out1: 3.06401  V
** sourceTransconductance: 3.39501  V


.END