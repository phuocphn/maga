** Name: two_stage_single_output_op_amp_40_9

.MACRO two_stage_single_output_op_amp_40_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=4e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=234e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=41e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=233e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=9e-6 W=20e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=63e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=20e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=41e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=234e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=24e-6
mSecondStage1StageBias13 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=233e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=20e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=343e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=9e-6 W=20e-6
mMainBias18 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=151e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_40_9

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 4.05501 mW
** Area: 10628 (mu_m)^2
** Transit frequency: 3.65401 MHz
** Transit frequency with error factor: 3.65006 MHz
** Slew rate: 5.61749 V/mu_s
** Phase margin: 60.7336°
** CMRR: 94 dB
** negPSRR: 104 dB
** posPSRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 1 V
** VcmMax: 3.53001 V
** VcmMin: 1.59001 V


** Expected Currents: 
** NormalTransistorNmos: 5.96491e+07 muA
** NormalTransistorPmos: -1.41916e+08 muA
** DiodeTransistorPmos: -1.26709e+07 muA
** NormalTransistorPmos: -1.26699e+07 muA
** NormalTransistorPmos: -1.26689e+07 muA
** DiodeTransistorPmos: -1.26699e+07 muA
** NormalTransistorNmos: 2.53391e+07 muA
** DiodeTransistorNmos: 2.53381e+07 muA
** NormalTransistorNmos: 1.26701e+07 muA
** NormalTransistorNmos: 1.26701e+07 muA
** NormalTransistorNmos: 5.74187e+08 muA
** DiodeTransistorNmos: 5.74188e+08 muA
** NormalTransistorPmos: -5.74186e+08 muA
** DiodeTransistorNmos: 1.41917e+08 muA
** NormalTransistorNmos: 1.41916e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.96499e+07 muA


** Expected Voltages: 
** ibias: 1.40201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.97601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.34801  V
** outSourceVoltageBiasXXnXX1: 0.674001  V
** outSourceVoltageBiasXXnXX2: 0.702001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.24801  V
** innerTransistorStack1Load1: 4.24901  V
** out1: 3.12201  V
** sourceTransconductance: 1.85001  V
** inner: 0.674001  V
** inner: 0.698001  V


.END