** Name: two_stage_single_output_op_amp_197_12

.MACRO two_stage_single_output_op_amp_197_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=2e-6 W=12e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=28e-6
mMainBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=7e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=426e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=371e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=157e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=168e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=426e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=12e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=157e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=375e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=79e-6
mSimpleFirstStageLoad19 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=129e-6
mSimpleFirstStageLoad20 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=129e-6
mSimpleFirstStageLoad21 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=180e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=577e-6
mMainBias23 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mSecondStage1Transconductor24 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad25 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=180e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.3001e-12
.EOM two_stage_single_output_op_amp_197_12

** Expected Performance Values: 
** Gain: 140 dB
** Power consumption: 10.4991 mW
** Area: 14990 (mu_m)^2
** Transit frequency: 9.47601 MHz
** Transit frequency with error factor: 9.4713 MHz
** Slew rate: 8.93071 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** VoutMax: 4.25 V
** VoutMin: 1.39001 V
** VcmMax: 4.84001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorNmos: 2.51761e+07 muA
** NormalTransistorPmos: -2.39719e+07 muA
** DiodeTransistorNmos: 1.58266e+08 muA
** DiodeTransistorNmos: 1.58265e+08 muA
** NormalTransistorNmos: 1.58264e+08 muA
** NormalTransistorNmos: 1.58265e+08 muA
** NormalTransistorPmos: -2.18071e+08 muA
** NormalTransistorPmos: -2.1807e+08 muA
** NormalTransistorPmos: -2.18069e+08 muA
** NormalTransistorPmos: -2.1807e+08 muA
** NormalTransistorNmos: 1.19612e+08 muA
** NormalTransistorNmos: 1.19611e+08 muA
** NormalTransistorNmos: 5.98061e+07 muA
** NormalTransistorNmos: 5.98061e+07 muA
** NormalTransistorNmos: 1.48267e+09 muA
** DiodeTransistorNmos: 1.48267e+09 muA
** NormalTransistorPmos: -1.48266e+09 muA
** NormalTransistorPmos: -1.48266e+09 muA
** DiodeTransistorNmos: 2.39711e+07 muA
** NormalTransistorNmos: 2.39701e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.21839e+08 muA
** DiodeTransistorPmos: -2.51769e+07 muA


** Expected Voltages: 
** ibias: 1.12001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.80001  V
** out: 2.5  V
** outFirstStage: 4.05601  V
** outSourceVoltageBiasXXnXX1: 0.900001  V
** outSourceVoltageBiasXXnXX2: 0.556001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.12801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.13901  V
** innerStageBias: 0.490001  V
** innerTransistorStack1Load2: 4.51001  V
** innerTransistorStack2Load1: 1.14001  V
** innerTransistorStack2Load2: 4.51001  V
** out1: 2.10501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.62001  V
** inner: 0.900001  V


.END