** Name: two_stage_single_output_op_amp_197_11

.MACRO two_stage_single_output_op_amp_197_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=39e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=57e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=5e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=110e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=146e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=26e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=39e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=45e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=10e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=599e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=127e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=57e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=45e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=423e-6
mMainBias16 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=201e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad19 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=442e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=366e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=599e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=442e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_197_11

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 9.59401 mW
** Area: 14144 (mu_m)^2
** Transit frequency: 3.83301 MHz
** Transit frequency with error factor: 3.8294 MHz
** Slew rate: 3.61239 V/mu_s
** Phase margin: 60.1606°
** CMRR: 128 dB
** VoutMax: 4.26001 V
** VoutMin: 0.890001 V
** VcmMax: 4.66001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 2.79218e+08 muA
** NormalTransistorNmos: 1.33415e+08 muA
** DiodeTransistorNmos: 5.39714e+08 muA
** DiodeTransistorNmos: 5.39713e+08 muA
** NormalTransistorNmos: 5.39714e+08 muA
** NormalTransistorNmos: 5.39713e+08 muA
** NormalTransistorPmos: -5.48284e+08 muA
** NormalTransistorPmos: -5.48283e+08 muA
** NormalTransistorPmos: -5.48284e+08 muA
** NormalTransistorPmos: -5.48283e+08 muA
** NormalTransistorNmos: 1.71411e+07 muA
** NormalTransistorNmos: 1.71401e+07 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 3.99652e+08 muA
** NormalTransistorNmos: 3.99651e+08 muA
** NormalTransistorPmos: -3.99651e+08 muA
** NormalTransistorPmos: -3.99652e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.79217e+08 muA
** DiodeTransistorPmos: -1.33414e+08 muA


** Expected Voltages: 
** ibias: 1.22801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.08501  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.21101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.10801  V
** innerStageBias: 0.576001  V
** innerTransistorStack1Load2: 4.77501  V
** innerTransistorStack2Load1: 1.10801  V
** innerTransistorStack2Load2: 4.77501  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.488001  V
** innerTransconductance: 4.63501  V


.END