** Name: two_stage_single_output_op_amp_26_5

.MACRO two_stage_single_output_op_amp_26_5 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=29e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=29e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=221e-6
mMainBias4 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=2e-6 W=10e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=286e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=256e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=539e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=29e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=279e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=29e-6
mMainBias11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=61e-6
mSimpleFirstStageTransconductor12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=155e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=256e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=286e-6
mMainBias15 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mSecondStage1StageBias16 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=539e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=155e-6
mMainBias18 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=168e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_26_5

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 4.14601 mW
** Area: 13577 (mu_m)^2
** Transit frequency: 4.13401 MHz
** Transit frequency with error factor: 4.13085 MHz
** Slew rate: 4.50335 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** negPSRR: 97 dB
** posPSRR: 99 dB
** VoutMax: 3.76001 V
** VoutMin: 0.460001 V
** VcmMax: 3.27001 V
** VcmMin: 0.610001 V


** Expected Currents: 
** NormalTransistorNmos: 4.72821e+07 muA
** NormalTransistorPmos: -1.71176e+08 muA
** DiodeTransistorNmos: 2.08111e+07 muA
** NormalTransistorNmos: 2.08101e+07 muA
** NormalTransistorNmos: 2.08111e+07 muA
** DiodeTransistorNmos: 2.08101e+07 muA
** NormalTransistorPmos: -4.1625e+07 muA
** DiodeTransistorPmos: -4.16259e+07 muA
** NormalTransistorPmos: -2.08119e+07 muA
** NormalTransistorPmos: -2.08119e+07 muA
** NormalTransistorNmos: 5.49196e+08 muA
** NormalTransistorPmos: -5.49195e+08 muA
** DiodeTransistorPmos: -5.49194e+08 muA
** DiodeTransistorNmos: 1.71177e+08 muA
** DiodeTransistorPmos: -4.72829e+07 muA
** NormalTransistorPmos: -4.72829e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.19701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.861001  V
** outInputVoltageBiasXXpXX1: 3.44401  V
** outSourceVoltageBiasXXpXX1: 4.22201  V
** outSourceVoltageBiasXXpXX2: 4.10001  V
** outVoltageBiasXXnXX0: 0.618001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.610001  V
** innerTransistorStack1Load1: 0.609001  V
** out1: 1.17401  V
** sourceTransconductance: 3.23701  V
** inner: 4.22201  V
** inner: 4.09401  V


.END