** Name: two_stage_single_output_op_amp_20_3

.MACRO two_stage_single_output_op_amp_20_3 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=126e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=11e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=4e-6 W=26e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=23e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=75e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=126e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=485e-6
mSimpleFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=46e-6
mMainBias11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=32e-6
mSimpleFirstStageTransconductor12 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=14e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=75e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=91e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSecondStage1StageBias16 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=4e-6 W=599e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=14e-6
mMainBias18 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=8e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_20_3

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 1.86901 mW
** Area: 7469 (mu_m)^2
** Transit frequency: 6.52101 MHz
** Transit frequency with error factor: 6.50939 MHz
** Slew rate: 9.33207 V/mu_s
** Phase margin: 63.5984°
** CMRR: 99 dB
** negPSRR: 100 dB
** posPSRR: 182 dB
** VoutMax: 3.39001 V
** VoutMin: 0.150001 V
** VcmMax: 3.05001 V
** VcmMin: 0.260001 V


** Expected Currents: 
** NormalTransistorNmos: 2.12021e+07 muA
** NormalTransistorPmos: -1.26909e+07 muA
** NormalTransistorPmos: -2.02489e+07 muA
** DiodeTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorPmos: -6.85709e+07 muA
** DiodeTransistorPmos: -6.85719e+07 muA
** NormalTransistorPmos: -3.42849e+07 muA
** NormalTransistorPmos: -3.42849e+07 muA
** NormalTransistorNmos: 2.30991e+08 muA
** NormalTransistorPmos: -2.3099e+08 muA
** NormalTransistorPmos: -2.30989e+08 muA
** DiodeTransistorNmos: 1.26901e+07 muA
** DiodeTransistorNmos: 2.02481e+07 muA
** DiodeTransistorPmos: -2.12029e+07 muA
** NormalTransistorPmos: -2.12039e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.82801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.41801  V
** outSourceVoltageBiasXXpXX1: 4.20901  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX0: 0.559001  V
** outVoltageBiasXXnXX1: 0.820001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.43301  V
** innerStageBias: 3.68501  V
** inner: 4.20801  V


.END