** Name: two_stage_single_output_op_amp_97_9

.MACRO two_stage_single_output_op_amp_97_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=561e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=9e-6
mTelescopicFirstStageLoad5 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=10e-6 W=18e-6
mMainBias7 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=11e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=32e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=43e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=43e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=561e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=32e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=26e-6
mTelescopicFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=206e-6
mTelescopicFirstStageLoad18 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=10e-6 W=18e-6
mMainBias19 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=89e-6
mMainBias20 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=20e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_97_9

** Expected Performance Values: 
** Gain: 131 dB
** Power consumption: 14.9991 mW
** Area: 3908 (mu_m)^2
** Transit frequency: 4.81301 MHz
** Transit frequency with error factor: 4.81319 MHz
** Slew rate: 7.05861 V/mu_s
** Phase margin: 69.9009°
** CMRR: 133 dB
** VoutMax: 4.11001 V
** VoutMin: 0.900001 V
** VcmMax: 3.39001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorNmos: 6.15501e+06 muA
** NormalTransistorPmos: -5.07189e+07 muA
** NormalTransistorPmos: -1.13839e+07 muA
** NormalTransistorNmos: 1.02391e+07 muA
** NormalTransistorNmos: 1.02391e+07 muA
** DiodeTransistorPmos: -1.02399e+07 muA
** NormalTransistorPmos: -1.02409e+07 muA
** NormalTransistorPmos: -1.02399e+07 muA
** DiodeTransistorPmos: -1.02409e+07 muA
** NormalTransistorNmos: 3.18601e+07 muA
** NormalTransistorNmos: 1.02381e+07 muA
** NormalTransistorNmos: 1.02381e+07 muA
** NormalTransistorNmos: 2.90116e+09 muA
** DiodeTransistorNmos: 2.90116e+09 muA
** NormalTransistorPmos: -2.90115e+09 muA
** DiodeTransistorNmos: 5.07201e+07 muA
** NormalTransistorNmos: 5.07201e+07 muA
** DiodeTransistorNmos: 1.13831e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.15599e+06 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.54401  V
** outInputVoltageBiasXXnXX1: 1.30201  V
** outSourceVoltageBiasXXnXX1: 0.651001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 3.93301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.25201  V
** innerTransistorStack2Load2: 4.25701  V
** out1: 3.12601  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.651001  V


.END