** Name: two_stage_single_output_op_amp_10_10

.MACRO two_stage_single_output_op_amp_10_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=146e-6
mMainBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mSimpleFirstStageTransconductor4 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=47e-6
mSimpleFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=113e-6
mSecondStage1StageBias6 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=473e-6
mSimpleFirstStageTransconductor7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=47e-6
mMainBias8 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=244e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=146e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=522e-6
mSecondStage1Transconductor11 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=316e-6
mSimpleFirstStageLoad12 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=60e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.6001e-12
.EOM two_stage_single_output_op_amp_10_10

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 5.16801 mW
** Area: 7140 (mu_m)^2
** Transit frequency: 3.61401 MHz
** Transit frequency with error factor: 3.60862 MHz
** Slew rate: 9.47903 V/mu_s
** Phase margin: 60.1606°
** CMRR: 95 dB
** negPSRR: 113 dB
** posPSRR: 93 dB
** VoutMax: 4.25 V
** VoutMin: 0.240001 V
** VcmMax: 4.30001 V
** VcmMin: 1.07001 V


** Expected Currents: 
** NormalTransistorNmos: 3.04602e+08 muA
** DiodeTransistorPmos: -6.93319e+07 muA
** NormalTransistorPmos: -6.93319e+07 muA
** NormalTransistorPmos: -6.93319e+07 muA
** NormalTransistorNmos: 1.38663e+08 muA
** NormalTransistorNmos: 6.93311e+07 muA
** NormalTransistorNmos: 6.93311e+07 muA
** NormalTransistorNmos: 5.80415e+08 muA
** NormalTransistorPmos: -5.80414e+08 muA
** NormalTransistorPmos: -5.80415e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.04601e+08 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.00501  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.15301  V
** innerTransistorStack2Load1: 4.50401  V
** sourceTransconductance: 1.67601  V
** innerTransconductance: 4.56901  V


.END