** Name: symmetrical_op_amp49

.MACRO symmetrical_op_amp49 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=22e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=62e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=43e-6
mSymmetricalFirstStageLoad4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=62e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=175e-6
mSymmetricalFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=117e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=36e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=62e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=62e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=7e-6 W=210e-6
mSecondStage1Transconductor12 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=7e-6 W=210e-6
mMainBias13 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=121e-6
mSymmetricalFirstStageStageBias14 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=117e-6
mSecondStage1StageBias15 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=175e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias17 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mSymmetricalFirstStageTransconductor18 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=104e-6
mMainBias19 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=129e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=146e-6
mSymmetricalFirstStageTransconductor21 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=104e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp49

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 3.89001 mW
** Area: 7329 (mu_m)^2
** Transit frequency: 5.26401 MHz
** Transit frequency with error factor: 5.26357 MHz
** Slew rate: 5.88146 V/mu_s
** Phase margin: 72.7657°
** CMRR: 154 dB
** negPSRR: 53 dB
** posPSRR: 89 dB
** VoutMax: 4.49001 V
** VoutMin: 0.300001 V
** VcmMax: 3.22001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 3.65522e+08 muA
** NormalTransistorPmos: -1.30789e+08 muA
** NormalTransistorPmos: -2.43329e+07 muA
** DiodeTransistorNmos: 5.93111e+07 muA
** DiodeTransistorNmos: 5.93111e+07 muA
** NormalTransistorPmos: -1.18623e+08 muA
** DiodeTransistorPmos: -1.18622e+08 muA
** NormalTransistorPmos: -5.93119e+07 muA
** NormalTransistorPmos: -5.93119e+07 muA
** NormalTransistorNmos: 5.90431e+07 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorPmos: -5.90439e+07 muA
** NormalTransistorPmos: -5.90449e+07 muA
** DiodeTransistorPmos: -5.96409e+07 muA
** NormalTransistorNmos: 5.96401e+07 muA
** NormalTransistorNmos: 5.96391e+07 muA
** DiodeTransistorNmos: 1.3079e+08 muA
** DiodeTransistorNmos: 2.43321e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -3.65521e+08 muA


** Expected Voltages: 
** ibias: 3.39601  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.708001  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 4.07101  V
** inputVoltageBiasXXnXX0: 0.732001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.24201  V
** innerStageBias: 4.40001  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V
** inner: 4.19601  V


.END