** Name: two_stage_single_output_op_amp_169_5

.MACRO two_stage_single_output_op_amp_169_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=10e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=7e-6 W=21e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=21e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=7e-6 W=7e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=19e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=470e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=10e-6
mSimpleFirstStageLoad9 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=36e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=42e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=42e-6
mMainBias12 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSecondStage1Transconductor13 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=545e-6
mSimpleFirstStageLoad14 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=36e-6
mMainBias15 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=59e-6
mSimpleFirstStageTransconductor16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=148e-6
mSimpleFirstStageStageBias17 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=44e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=21e-6
mSimpleFirstStageStageBias19 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=7e-6 W=214e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=470e-6
mSimpleFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=7e-6 W=21e-6
mSimpleFirstStageTransconductor23 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=148e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_169_5

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 7.90601 mW
** Area: 8656 (mu_m)^2
** Transit frequency: 4.45801 MHz
** Transit frequency with error factor: 4.45678 MHz
** Slew rate: 4.7226 V/mu_s
** Phase margin: 60.1606°
** CMRR: 100 dB
** VoutMax: 3.27001 V
** VoutMin: 0.310001 V
** VcmMax: 3.07001 V
** VcmMin: -0.25 V


** Expected Currents: 
** NormalTransistorNmos: 5.81021e+07 muA
** NormalTransistorNmos: 4.96901e+06 muA
** DiodeTransistorPmos: -3.04599e+07 muA
** DiodeTransistorPmos: -3.04599e+07 muA
** NormalTransistorPmos: -3.04599e+07 muA
** NormalTransistorPmos: -3.04599e+07 muA
** NormalTransistorNmos: 4.12001e+07 muA
** NormalTransistorNmos: 4.12011e+07 muA
** NormalTransistorNmos: 4.12001e+07 muA
** NormalTransistorNmos: 4.12011e+07 muA
** NormalTransistorPmos: -2.14829e+07 muA
** NormalTransistorPmos: -2.14839e+07 muA
** NormalTransistorPmos: -1.07409e+07 muA
** NormalTransistorPmos: -1.07409e+07 muA
** NormalTransistorNmos: 1.42569e+09 muA
** NormalTransistorPmos: -1.42568e+09 muA
** DiodeTransistorPmos: -1.42568e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.81029e+07 muA
** NormalTransistorPmos: -5.81039e+07 muA
** DiodeTransistorPmos: -4.96999e+06 muA
** DiodeTransistorPmos: -4.96899e+06 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.90301  V
** out: 2.5  V
** outFirstStage: 0.711001  V
** outInputVoltageBiasXXpXX1: 2.70201  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 3.85101  V
** outSourceVoltageBiasXXpXX2: 3.99701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerSourceLoad1: 3.68601  V
** innerStageBias: 3.66501  V
** innerTransistorStack1Load2: 0.546001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.546001  V
** sourceTransconductance: 3.23201  V
** inner: 3.84901  V


.END