** Name: two_stage_single_output_op_amp_59_5

.MACRO two_stage_single_output_op_amp_59_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=16e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=80e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=7e-6 W=23e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=6e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=379e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
mMainBias11 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=15e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=10e-6 W=244e-6
mFoldedCascodeFirstStageLoad13 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=26e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=25e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=37e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=80e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=198e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=198e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=7e-6 W=206e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=6e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=379e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=8e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.80001e-12
.EOM two_stage_single_output_op_amp_59_5

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 3.44701 mW
** Area: 12242 (mu_m)^2
** Transit frequency: 4.29401 MHz
** Transit frequency with error factor: 4.29358 MHz
** Slew rate: 4.34426 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** VoutMax: 3.40001 V
** VoutMin: 0.540001 V
** VcmMax: 3.03001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 9.61901e+06 muA
** NormalTransistorNmos: 5.77101e+06 muA
** NormalTransistorNmos: 2.09031e+07 muA
** NormalTransistorNmos: 3.16171e+07 muA
** NormalTransistorNmos: 2.09031e+07 muA
** NormalTransistorNmos: 3.16171e+07 muA
** NormalTransistorPmos: -2.09039e+07 muA
** NormalTransistorPmos: -2.09039e+07 muA
** DiodeTransistorPmos: -2.09039e+07 muA
** NormalTransistorPmos: -2.14309e+07 muA
** NormalTransistorPmos: -2.14319e+07 muA
** NormalTransistorPmos: -1.07149e+07 muA
** NormalTransistorPmos: -1.07149e+07 muA
** NormalTransistorNmos: 6.00752e+08 muA
** NormalTransistorPmos: -6.00751e+08 muA
** DiodeTransistorPmos: -6.00752e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.61999e+06 muA
** NormalTransistorPmos: -9.62099e+06 muA
** DiodeTransistorPmos: -5.77199e+06 muA
** DiodeTransistorPmos: -5.77299e+06 muA


** Expected Voltages: 
** ibias: 1.15201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.08001  V
** out: 2.5  V
** outFirstStage: 0.947001  V
** outInputVoltageBiasXXpXX1: 2.83601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.91801  V
** outSourceVoltageBiasXXpXX2: 3.95901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.22601  V
** innerStageBias: 3.84501  V
** out1: 3.11901  V
** sourceGCC1: 0.528001  V
** sourceGCC2: 0.528001  V
** sourceTransconductance: 3.22901  V
** inner: 3.91701  V


.END