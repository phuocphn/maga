** Name: two_stage_single_output_op_amp_57_11

.MACRO two_stage_single_output_op_amp_57_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=6e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=151e-6
mSecondStage1StageBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=59e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=190e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=16e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=75e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=75e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=563e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=150e-6
mSecondStage1StageBias11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=123e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=16e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=53e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=10e-6 W=181e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=40e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=40e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=6e-6 W=221e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=584e-6
mSecondStage1Transconductor19 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=6e-6 W=532e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=151e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.70001e-12
.EOM two_stage_single_output_op_amp_57_11

** Expected Performance Values: 
** Gain: 132 dB
** Power consumption: 3.07201 mW
** Area: 14998 (mu_m)^2
** Transit frequency: 2.79301 MHz
** Transit frequency with error factor: 2.78944 MHz
** Slew rate: 3.72707 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** VoutMax: 4.25 V
** VoutMin: 0.890001 V
** VcmMax: 3.12001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 9.98401e+07 muA
** NormalTransistorNmos: 3.46621e+07 muA
** NormalTransistorNmos: 3.25871e+07 muA
** NormalTransistorNmos: 4.90491e+07 muA
** NormalTransistorNmos: 3.25871e+07 muA
** NormalTransistorNmos: 4.90491e+07 muA
** DiodeTransistorPmos: -3.25879e+07 muA
** NormalTransistorPmos: -3.25879e+07 muA
** NormalTransistorPmos: -3.29269e+07 muA
** NormalTransistorPmos: -3.29279e+07 muA
** NormalTransistorPmos: -1.64629e+07 muA
** NormalTransistorPmos: -1.64629e+07 muA
** NormalTransistorNmos: 3.71829e+08 muA
** NormalTransistorNmos: 3.71828e+08 muA
** NormalTransistorPmos: -3.71828e+08 muA
** NormalTransistorPmos: -3.71829e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.98409e+07 muA
** DiodeTransistorPmos: -3.46629e+07 muA


** Expected Voltages: 
** ibias: 1.20501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.16801  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX2: 4.11601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.47301  V
** out1: 4.16601  V
** sourceGCC1: 0.530001  V
** sourceGCC2: 0.530001  V
** sourceTransconductance: 3.27801  V
** innerStageBias: 0.472001  V
** innerTransconductance: 4.73201  V


.END