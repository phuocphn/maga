** Name: two_stage_single_output_op_amp_80_12

.MACRO two_stage_single_output_op_amp_80_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=52e-6
mMainBias2 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=13e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=45e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=510e-6
mMainBias6 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=6e-6
mMainBias7 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=63e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=108e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=63e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=63e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=115e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=115e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=45e-6
mMainBias15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mMainBias16 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=52e-6
mSecondStage1StageBias17 out inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=510e-6
mFoldedCascodeFirstStageLoad18 outFirstStage inputVoltageBiasXXnXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=108e-6
mMainBias19 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=20e-6
mFoldedCascodeFirstStageLoad20 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=298e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=566e-6
mFoldedCascodeFirstStageLoad22 FirstStageYsourceGCC2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=566e-6
mSecondStage1Transconductor23 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=347e-6
mMainBias24 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=510e-6
mMainBias25 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=345e-6
mSecondStage1Transconductor26 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=599e-6
mFoldedCascodeFirstStageLoad27 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=298e-6
mMainBias28 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=114e-6
mMainBias29 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=46e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.1001e-12
.EOM two_stage_single_output_op_amp_80_12

** Expected Performance Values: 
** Gain: 176 dB
** Power consumption: 6.02501 mW
** Area: 14985 (mu_m)^2
** Transit frequency: 3.85701 MHz
** Transit frequency with error factor: 3.85745 MHz
** Slew rate: 3.50334 V/mu_s
** Phase margin: 60.1606°
** CMRR: 149 dB
** VoutMax: 4.25 V
** VoutMin: 0.790001 V
** VcmMax: 5.24001 V
** VcmMin: 1.47001 V


** Expected Currents: 
** NormalTransistorNmos: 2.53041e+07 muA
** NormalTransistorPmos: -7.44399e+06 muA
** NormalTransistorPmos: -1.82129e+07 muA
** NormalTransistorPmos: -8.20129e+07 muA
** NormalTransistorPmos: -5.49279e+07 muA
** NormalTransistorPmos: -6.03049e+07 muA
** NormalTransistorPmos: -9.15949e+07 muA
** NormalTransistorPmos: -6.03049e+07 muA
** NormalTransistorPmos: -9.15949e+07 muA
** NormalTransistorNmos: 6.03041e+07 muA
** NormalTransistorNmos: 6.03031e+07 muA
** NormalTransistorNmos: 6.03041e+07 muA
** NormalTransistorNmos: 6.03031e+07 muA
** NormalTransistorNmos: 6.25811e+07 muA
** DiodeTransistorNmos: 6.25801e+07 muA
** NormalTransistorNmos: 3.12911e+07 muA
** NormalTransistorNmos: 3.12911e+07 muA
** NormalTransistorNmos: 8.13859e+08 muA
** DiodeTransistorNmos: 8.13858e+08 muA
** NormalTransistorPmos: -8.13858e+08 muA
** NormalTransistorPmos: -8.13859e+08 muA
** DiodeTransistorNmos: 7.44301e+06 muA
** DiodeTransistorNmos: 1.82121e+07 muA
** NormalTransistorNmos: 1.82111e+07 muA
** DiodeTransistorNmos: 8.20121e+07 muA
** NormalTransistorNmos: 8.20131e+07 muA
** DiodeTransistorNmos: 5.49271e+07 muA
** DiodeTransistorPmos: -2.53049e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.19801  V
** inputVoltageBiasXXnXX3: 0.917001  V
** out: 2.5  V
** outFirstStage: 4.07401  V
** outInputVoltageBiasXXnXX1: 1.32201  V
** outSourceVoltageBiasXXnXX1: 0.661001  V
** outSourceVoltageBiasXXnXX2: 0.599001  V
** outVoltageBiasXXnXX0: 0.677001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.63801  V
** inner: 0.659001  V
** inner: 0.600001  V


.END