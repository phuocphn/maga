** Name: two_stage_single_output_op_amp_65_11

.MACRO two_stage_single_output_op_amp_65_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=8e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=436e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=84e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=209e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=209e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=500e-6
mMainBias9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=325e-6
mSecondStage1StageBias10 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=356e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=84e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=113e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=541e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=195e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=195e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=74e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=127e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=127e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=340e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=186e-6
mSecondStage1Transconductor21 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=207e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=74e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.7001e-12
.EOM two_stage_single_output_op_amp_65_11

** Expected Performance Values: 
** Gain: 163 dB
** Power consumption: 6.75401 mW
** Area: 9593 (mu_m)^2
** Transit frequency: 2.69101 MHz
** Transit frequency with error factor: 2.69121 MHz
** Slew rate: 9.26965 V/mu_s
** Phase margin: 64.7443°
** CMRR: 132 dB
** VoutMax: 4.25 V
** VoutMin: 0.740001 V
** VcmMax: 3.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.24909e+08 muA
** NormalTransistorNmos: 1.10852e+08 muA
** NormalTransistorNmos: 1.36613e+08 muA
** NormalTransistorNmos: 2.05026e+08 muA
** NormalTransistorNmos: 1.36613e+08 muA
** NormalTransistorNmos: 2.05026e+08 muA
** NormalTransistorPmos: -1.36612e+08 muA
** NormalTransistorPmos: -1.36613e+08 muA
** NormalTransistorPmos: -1.36612e+08 muA
** NormalTransistorPmos: -1.36613e+08 muA
** NormalTransistorPmos: -1.36828e+08 muA
** NormalTransistorPmos: -1.36829e+08 muA
** NormalTransistorPmos: -6.84139e+07 muA
** NormalTransistorPmos: -6.84139e+07 muA
** NormalTransistorNmos: 4.95065e+08 muA
** NormalTransistorNmos: 4.95064e+08 muA
** NormalTransistorPmos: -4.95064e+08 muA
** NormalTransistorPmos: -4.95065e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.24908e+08 muA
** DiodeTransistorPmos: -1.10851e+08 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.05001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX2: 4.26701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40001  V
** innerTransistorStack1Load2: 4.57001  V
** innerTransistorStack2Load2: 4.57001  V
** out1: 4.23801  V
** sourceGCC1: 0.532001  V
** sourceGCC2: 0.532001  V
** sourceTransconductance: 3.61101  V
** innerStageBias: 0.547001  V
** innerTransconductance: 4.61401  V


.END