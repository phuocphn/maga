** Name: two_stage_single_output_op_amp_144_10

.MACRO two_stage_single_output_op_amp_144_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=242e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=45e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=151e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=35e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=242e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=41e-6
mMainBias8 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=107e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=563e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=73e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=35e-6
mMainBias12 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=134e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=591e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=591e-6
mSimpleFirstStageLoad15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=536e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=567e-6
mSecondStage1Transconductor17 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=600e-6
mSimpleFirstStageLoad18 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=536e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.40001e-12
.EOM two_stage_single_output_op_amp_144_10

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 13.0411 mW
** Area: 14538 (mu_m)^2
** Transit frequency: 7.07701 MHz
** Transit frequency with error factor: 7.0726 MHz
** Slew rate: 7.58524 V/mu_s
** Phase margin: 60.1606°
** CMRR: 119 dB
** VoutMax: 4.25 V
** VoutMin: 0.220001 V
** VcmMax: 4.66001 V
** VcmMin: 0.800001 V


** Expected Currents: 
** NormalTransistorNmos: 1.52301e+08 muA
** NormalTransistorNmos: 1.89965e+08 muA
** NormalTransistorNmos: 7.02212e+08 muA
** NormalTransistorNmos: 7.02211e+08 muA
** DiodeTransistorNmos: 7.02212e+08 muA
** NormalTransistorPmos: -7.30948e+08 muA
** NormalTransistorPmos: -7.30948e+08 muA
** NormalTransistorPmos: -7.30947e+08 muA
** NormalTransistorPmos: -7.30948e+08 muA
** NormalTransistorNmos: 5.74741e+07 muA
** NormalTransistorNmos: 2.87371e+07 muA
** NormalTransistorNmos: 2.87371e+07 muA
** NormalTransistorNmos: 7.94081e+08 muA
** NormalTransistorPmos: -7.9408e+08 muA
** NormalTransistorPmos: -7.94081e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.523e+08 muA
** DiodeTransistorPmos: -1.89964e+08 muA


** Expected Voltages: 
** ibias: 0.629001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.15501  V
** outVoltageBiasXXpXX2: 4.17201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.958001  V
** innerTransistorStack1Load2: 4.72701  V
** innerTransistorStack2Load2: 4.72701  V
** out1: 2.11301  V
** sourceTransconductance: 1.92401  V
** innerTransconductance: 4.71901  V


.END