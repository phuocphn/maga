** Name: two_stage_single_output_op_amp_43_6

.MACRO two_stage_single_output_op_amp_43_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=54e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=157e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=9e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=470e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=138e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=322e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=322e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=569e-6
mSecondStage1Transconductor11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=389e-6
mFoldedCascodeFirstStageLoad12 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=138e-6
mMainBias13 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=98e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=98e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=494e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
mMainBias18 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=102e-6
mSecondStage1StageBias19 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=470e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=157e-6
mMainBias21 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=85e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11e-12
.EOM two_stage_single_output_op_amp_43_6

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 12.2381 mW
** Area: 8827 (mu_m)^2
** Transit frequency: 9.47901 MHz
** Transit frequency with error factor: 9.44308 MHz
** Slew rate: 31.8447 V/mu_s
** Phase margin: 60.1606°
** CMRR: 85 dB
** VoutMax: 3.46001 V
** VoutMin: 0.550001 V
** VcmMax: 3.35001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorPmos: -8.55959e+07 muA
** NormalTransistorPmos: -1.0285e+08 muA
** NormalTransistorNmos: 3.64532e+08 muA
** NormalTransistorNmos: 6.13291e+08 muA
** NormalTransistorNmos: 3.64532e+08 muA
** NormalTransistorNmos: 6.13291e+08 muA
** DiodeTransistorPmos: -3.64531e+08 muA
** NormalTransistorPmos: -3.64531e+08 muA
** NormalTransistorPmos: -4.97516e+08 muA
** NormalTransistorPmos: -2.48757e+08 muA
** NormalTransistorPmos: -2.48757e+08 muA
** NormalTransistorNmos: 9.9352e+08 muA
** NormalTransistorNmos: 9.93521e+08 muA
** NormalTransistorPmos: -9.93519e+08 muA
** DiodeTransistorPmos: -9.9352e+08 muA
** DiodeTransistorNmos: 8.55951e+07 muA
** DiodeTransistorNmos: 1.02851e+08 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90489e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.10001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.655001  V
** outInputVoltageBiasXXpXX1: 2.89601  V
** outSourceVoltageBiasXXpXX1: 3.94801  V
** outVoltageBiasXXnXX1: 1.06001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.07401  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.81401  V
** innerTransconductance: 0.353001  V
** inner: 3.94501  V


.END