** Name: two_stage_single_output_op_amp_77_10

.MACRO two_stage_single_output_op_amp_77_10 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=374e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=4e-6 W=350e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mMainBias4 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=27e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=442e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=208e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=4e-6 W=350e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=17e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=119e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=374e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=82e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=242e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerOutputLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=277e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=564e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=564e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=371e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=599e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=277e-6
mMainBias22 outVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=588e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.1001e-12
.EOM two_stage_single_output_op_amp_77_10

** Expected Performance Values: 
** Gain: 115 dB
** Power consumption: 10.3901 mW
** Area: 14513 (mu_m)^2
** Transit frequency: 4.02001 MHz
** Transit frequency with error factor: 4.01953 MHz
** Slew rate: 18.3217 V/mu_s
** Phase margin: 60.1606°
** CMRR: 127 dB
** VoutMax: 4.25 V
** VoutMin: 0.160001 V
** VcmMax: 5.22001 V
** VcmMin: 1.87001 V


** Expected Currents: 
** NormalTransistorNmos: 9.13791e+07 muA
** NormalTransistorNmos: 2.67186e+08 muA
** NormalTransistorPmos: -3.55441e+08 muA
** NormalTransistorPmos: -2.2448e+08 muA
** NormalTransistorPmos: -3.40933e+08 muA
** NormalTransistorPmos: -2.2448e+08 muA
** NormalTransistorPmos: -3.40933e+08 muA
** DiodeTransistorNmos: 2.24481e+08 muA
** DiodeTransistorNmos: 2.2448e+08 muA
** NormalTransistorNmos: 2.24481e+08 muA
** NormalTransistorNmos: 2.2448e+08 muA
** NormalTransistorNmos: 2.32904e+08 muA
** NormalTransistorNmos: 2.32903e+08 muA
** NormalTransistorNmos: 1.16453e+08 muA
** NormalTransistorNmos: 1.16453e+08 muA
** NormalTransistorNmos: 6.72078e+08 muA
** NormalTransistorPmos: -6.72077e+08 muA
** NormalTransistorPmos: -6.72078e+08 muA
** DiodeTransistorNmos: 3.55442e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.13799e+07 muA
** DiodeTransistorPmos: -2.67185e+08 muA


** Expected Voltages: 
** ibias: 0.567001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.11801  V
** outVoltageBiasXXnXX1: 0.971001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.25301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.15201  V
** innerStageBias: 0.414001  V
** innerTransistorStack1Load2: 0.579001  V
** innerTransistorStack2Load2: 0.578001  V
** sourceGCC1: 4.61701  V
** sourceGCC2: 4.61701  V
** sourceTransconductance: 1.34501  V
** innerTransconductance: 4.68201  V


.END