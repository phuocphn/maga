** Name: two_stage_single_output_op_amp_189_8

.MACRO two_stage_single_output_op_amp_189_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=37e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=9e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=285e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=87e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=20e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=12e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=37e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=21e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=476e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=318e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=22e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=12e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=323e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=323e-6
mSimpleFirstStageLoad17 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=592e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=368e-6
mSimpleFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=592e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_189_8

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 4.49901 mW
** Area: 12334 (mu_m)^2
** Transit frequency: 2.58901 MHz
** Transit frequency with error factor: 2.58597 MHz
** Slew rate: 4.27044 V/mu_s
** Phase margin: 63.0254°
** CMRR: 117 dB
** VoutMax: 4.25 V
** VoutMin: 0.740001 V
** VcmMax: 4.86001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 5.09541e+07 muA
** NormalTransistorNmos: 1.7592e+08 muA
** NormalTransistorNmos: 1.75921e+08 muA
** DiodeTransistorNmos: 1.7592e+08 muA
** NormalTransistorPmos: -1.85918e+08 muA
** NormalTransistorPmos: -1.85919e+08 muA
** NormalTransistorPmos: -1.85919e+08 muA
** NormalTransistorPmos: -1.85919e+08 muA
** NormalTransistorNmos: 1.99991e+07 muA
** NormalTransistorNmos: 1.99981e+07 muA
** NormalTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 4.67056e+08 muA
** NormalTransistorNmos: 4.67055e+08 muA
** NormalTransistorPmos: -4.67055e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.09549e+07 muA
** DiodeTransistorPmos: -5.09559e+07 muA


** Expected Voltages: 
** ibias: 1.125  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.38601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.12401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.570001  V
** innerTransistorStack1Load2: 4.17901  V
** innerTransistorStack2Load2: 4.17901  V
** out1: 2.09501  V
** sourceTransconductance: 1.83201  V
** innerStageBias: 0.533001  V


.END