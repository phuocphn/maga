** Name: two_stage_single_output_op_amp_64_4

.MACRO two_stage_single_output_op_amp_64_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=146e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=25e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=58e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=6e-6 W=120e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=9e-6 W=102e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=231e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=23e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=88e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=88e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=104e-6
mSecondStage1Transconductor13 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageLoad14 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=23e-6
mMainBias15 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=27e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=57e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=57e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=9e-6 W=231e-6
mSecondStage1StageBias20 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=59e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=102e-6
mMainBias22 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=33e-6
mSecondStage1StageBias23 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=6e-6 W=599e-6
mFoldedCascodeFirstStageLoad24 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=58e-6
mMainBias25 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=156e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.30001e-12
.EOM two_stage_single_output_op_amp_64_4

** Expected Performance Values: 
** Gain: 183 dB
** Power consumption: 2.58601 mW
** Area: 14997 (mu_m)^2
** Transit frequency: 2.66601 MHz
** Transit frequency with error factor: 2.66631 MHz
** Slew rate: 3.92229 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 3.45001 V
** VoutMin: 0.370001 V
** VcmMax: 3.16001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.02851e+07 muA
** NormalTransistorPmos: -2.63987e+08 muA
** NormalTransistorPmos: -5.58089e+07 muA
** NormalTransistorNmos: 2.19041e+07 muA
** NormalTransistorNmos: 3.36021e+07 muA
** NormalTransistorNmos: 2.19041e+07 muA
** NormalTransistorNmos: 3.36021e+07 muA
** DiodeTransistorPmos: -2.19049e+07 muA
** DiodeTransistorPmos: -2.19059e+07 muA
** NormalTransistorPmos: -2.19049e+07 muA
** NormalTransistorPmos: -2.19059e+07 muA
** NormalTransistorPmos: -2.33989e+07 muA
** DiodeTransistorPmos: -2.33999e+07 muA
** NormalTransistorPmos: -1.16989e+07 muA
** NormalTransistorPmos: -1.16989e+07 muA
** NormalTransistorNmos: 9.98411e+07 muA
** NormalTransistorNmos: 9.98401e+07 muA
** NormalTransistorPmos: -9.98419e+07 muA
** NormalTransistorPmos: -9.98409e+07 muA
** DiodeTransistorNmos: 2.63988e+08 muA
** DiodeTransistorNmos: 5.58081e+07 muA
** DiodeTransistorPmos: -1.02859e+07 muA
** NormalTransistorPmos: -1.02869e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.95401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.42001  V
** outSourceVoltageBiasXXpXX1: 4.21001  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX1: 0.905001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.03001  V
** innerTransistorStack2Load2: 4.02901  V
** out1: 3.26001  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.32601  V
** innerStageBias: 3.75401  V
** innerTransconductance: 0.275001  V
** inner: 4.20901  V


.END