** Name: two_stage_single_output_op_amp_58_7

.MACRO two_stage_single_output_op_amp_58_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=149e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=178e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=120e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=109e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=85e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=85e-6
mSecondStage1StageBias9 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=599e-6
mFoldedCascodeFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=109e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=257e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=257e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=120e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=178e-6
mMainBias17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=136e-6
mMainBias18 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=320e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.8001e-12
.EOM two_stage_single_output_op_amp_58_7

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 10.7661 mW
** Area: 5506 (mu_m)^2
** Transit frequency: 10.0501 MHz
** Transit frequency with error factor: 10.0377 MHz
** Slew rate: 10.2169 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** VoutMax: 4.65001 V
** VoutMin: 0.160001 V
** VcmMax: 3.03001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorPmos: -1.38571e+08 muA
** NormalTransistorPmos: -3.19693e+08 muA
** NormalTransistorNmos: 1.2124e+08 muA
** NormalTransistorNmos: 1.82376e+08 muA
** NormalTransistorNmos: 1.2124e+08 muA
** NormalTransistorNmos: 1.82376e+08 muA
** DiodeTransistorPmos: -1.21239e+08 muA
** NormalTransistorPmos: -1.21239e+08 muA
** NormalTransistorPmos: -1.22269e+08 muA
** DiodeTransistorPmos: -1.22268e+08 muA
** NormalTransistorPmos: -6.11349e+07 muA
** NormalTransistorPmos: -6.11349e+07 muA
** NormalTransistorNmos: 1.31024e+09 muA
** NormalTransistorPmos: -1.31023e+09 muA
** DiodeTransistorNmos: 1.38572e+08 muA
** DiodeTransistorNmos: 3.19694e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.19701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.08501  V
** outSourceVoltageBiasXXpXX1: 4.10001  V
** outVoltageBiasXXnXX1: 0.927001  V
** outVoltageBiasXXnXX2: 0.565001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.09701  V
** sourceGCC1: 0.360001  V
** sourceGCC2: 0.360001  V
** sourceTransconductance: 3.22701  V
** inner: 4.09401  V


.END