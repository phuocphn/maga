** Name: two_stage_single_output_op_amp_60_6

.MACRO two_stage_single_output_op_amp_60_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=9e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=115e-6
mMainBias4 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=4e-6 W=47e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=14e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=123e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=543e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=30e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=76e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=76e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=555e-6
mSecondStage1Transconductor12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=62e-6
mFoldedCascodeFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=30e-6
mMainBias14 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=6e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=115e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=46e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=46e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=123e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=14e-6
mMainBias20 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=47e-6
mSecondStage1StageBias21 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=4e-6 W=543e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=5e-6 W=117e-6
mMainBias23 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=133e-6
mMainBias24 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=16e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.80001e-12
.EOM two_stage_single_output_op_amp_60_6

** Expected Performance Values: 
** Gain: 184 dB
** Power consumption: 1.14901 mW
** Area: 14997 (mu_m)^2
** Transit frequency: 2.98601 MHz
** Transit frequency with error factor: 2.98622 MHz
** Slew rate: 3.94098 V/mu_s
** Phase margin: 60.1606°
** CMRR: 142 dB
** VoutMax: 4 V
** VoutMin: 0.410001 V
** VcmMax: 3.22001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.28601e+06 muA
** NormalTransistorPmos: -2.85019e+07 muA
** NormalTransistorPmos: -3.42999e+06 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 2.90501e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 2.90501e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -2.00089e+07 muA
** DiodeTransistorPmos: -2.00099e+07 muA
** NormalTransistorPmos: -1.00039e+07 muA
** NormalTransistorPmos: -1.00039e+07 muA
** NormalTransistorNmos: 1.17522e+08 muA
** NormalTransistorNmos: 1.17521e+08 muA
** NormalTransistorPmos: -1.17521e+08 muA
** DiodeTransistorPmos: -1.1752e+08 muA
** DiodeTransistorNmos: 2.85011e+07 muA
** DiodeTransistorNmos: 3.42901e+06 muA
** DiodeTransistorPmos: -2.28699e+06 muA
** NormalTransistorPmos: -2.28799e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.43201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.44401  V
** outSourceVoltageBiasXXpXX1: 4.22201  V
** outSourceVoltageBiasXXpXX2: 4.21701  V
** outVoltageBiasXXnXX1: 0.905001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.22001  V
** out1: 3.44201  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.28401  V
** innerTransconductance: 0.240001  V
** inner: 4.22101  V
** inner: 4.21401  V


.END