** Name: two_stage_single_output_op_amp_39_12

.MACRO two_stage_single_output_op_amp_39_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=32e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=8e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=81e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=231e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=5e-6 W=231e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=15e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=376e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=81e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=168e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias13 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=22e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=81e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=81e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=445e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=231e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=334e-6
mMainBias19 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=263e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=231e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.3001e-12
.EOM two_stage_single_output_op_amp_39_12

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 7.25001 mW
** Area: 14799 (mu_m)^2
** Transit frequency: 5.62701 MHz
** Transit frequency with error factor: 5.62429 MHz
** Slew rate: 5.30333 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** negPSRR: 116 dB
** posPSRR: 102 dB
** VoutMax: 4.25 V
** VoutMin: 1.53001 V
** VcmMax: 3.87001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 6.12701e+06 muA
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorPmos: -1.0702e+08 muA
** DiodeTransistorPmos: -5.14259e+07 muA
** NormalTransistorPmos: -5.14269e+07 muA
** NormalTransistorPmos: -5.14259e+07 muA
** DiodeTransistorPmos: -5.14269e+07 muA
** NormalTransistorNmos: 1.0285e+08 muA
** NormalTransistorNmos: 1.02849e+08 muA
** NormalTransistorNmos: 5.14251e+07 muA
** NormalTransistorNmos: 5.14251e+07 muA
** NormalTransistorNmos: 1.10211e+09 muA
** DiodeTransistorNmos: 1.10211e+09 muA
** NormalTransistorPmos: -1.1021e+09 muA
** NormalTransistorPmos: -1.1021e+09 muA
** DiodeTransistorNmos: 1.07021e+08 muA
** NormalTransistorNmos: 1.07021e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -6.12799e+06 muA
** DiodeTransistorPmos: -1.21839e+08 muA


** Expected Voltages: 
** ibias: 1.12101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.94001  V
** inputVoltageBiasXXpXX0: 4.00801  V
** out: 2.5  V
** outFirstStage: 4.00501  V
** outSourceVoltageBiasXXnXX1: 0.970001  V
** outSourceVoltageBiasXXnXX2: 0.556001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.27801  V
** innerStageBias: 0.490001  V
** innerTransistorStack1Load1: 4.27701  V
** out1: 3.46401  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.56901  V
** inner: 0.970001  V


.END