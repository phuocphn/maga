** Name: two_stage_single_output_op_amp_29_12

.MACRO two_stage_single_output_op_amp_29_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=5e-6 W=9e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=21e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=237e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=194e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=16e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=23e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=113e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=21e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=15e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=237e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=23e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=291e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=548e-6
mSecondStage1Transconductor17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=554e-6
mSimpleFirstStageLoad18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=194e-6
mMainBias19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=91e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.20001e-12
.EOM two_stage_single_output_op_amp_29_12

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 3.76401 mW
** Area: 12230 (mu_m)^2
** Transit frequency: 6.46101 MHz
** Transit frequency with error factor: 6.42494 MHz
** Slew rate: 12.7674 V/mu_s
** Phase margin: 60.1606°
** CMRR: 88 dB
** negPSRR: 114 dB
** posPSRR: 86 dB
** VoutMax: 4.62001 V
** VoutMin: 1.16001 V
** VcmMax: 4.66001 V
** VcmMin: 2 V


** Expected Currents: 
** NormalTransistorNmos: 5.74001e+06 muA
** NormalTransistorNmos: 1.11687e+08 muA
** NormalTransistorPmos: -3.22419e+07 muA
** DiodeTransistorPmos: -1.15432e+08 muA
** NormalTransistorPmos: -1.15432e+08 muA
** NormalTransistorNmos: 2.30864e+08 muA
** NormalTransistorNmos: 2.30863e+08 muA
** NormalTransistorNmos: 1.15433e+08 muA
** NormalTransistorNmos: 1.15433e+08 muA
** NormalTransistorNmos: 3.62299e+08 muA
** DiodeTransistorNmos: 3.62298e+08 muA
** NormalTransistorPmos: -3.62298e+08 muA
** NormalTransistorPmos: -3.62297e+08 muA
** DiodeTransistorNmos: 3.22411e+07 muA
** NormalTransistorNmos: 3.22401e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.74099e+06 muA
** DiodeTransistorPmos: -1.11686e+08 muA


** Expected Voltages: 
** ibias: 1.21501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.01201  V
** out: 2.5  V
** outFirstStage: 4.24301  V
** outInputVoltageBiasXXnXX1: 1.56801  V
** outSourceVoltageBiasXXnXX1: 0.784001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.462001  V
** out1: 4.25301  V
** sourceTransconductance: 1.40301  V
** innerTransconductance: 4.44101  V
** inner: 0.781001  V


.END