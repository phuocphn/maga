** Name: two_stage_single_output_op_amp_32_12

.MACRO two_stage_single_output_op_amp_32_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=6e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=166e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=33e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=412e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=149e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=63e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=149e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=123e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=33e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=166e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=42e-6
mSecondStage1StageBias13 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=412e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=123e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=459e-6
mSimpleFirstStageLoad16 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=149e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=349e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=467e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=9e-6 W=419e-6
mMainBias20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=212e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7e-12
.EOM two_stage_single_output_op_amp_32_12

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 8.94501 mW
** Area: 14859 (mu_m)^2
** Transit frequency: 6.93401 MHz
** Transit frequency with error factor: 6.93086 MHz
** Slew rate: 6.53547 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** negPSRR: 106 dB
** posPSRR: 100 dB
** VoutMax: 4.27001 V
** VoutMin: 0.890001 V
** VcmMax: 4.51001 V
** VcmMin: 1.48001 V


** Expected Currents: 
** NormalTransistorNmos: 7.00491e+07 muA
** NormalTransistorNmos: 7.56428e+08 muA
** NormalTransistorPmos: -2.31523e+08 muA
** NormalTransistorPmos: -2.34279e+07 muA
** NormalTransistorPmos: -2.34279e+07 muA
** DiodeTransistorPmos: -2.34279e+07 muA
** NormalTransistorNmos: 4.68531e+07 muA
** DiodeTransistorNmos: 4.68521e+07 muA
** NormalTransistorNmos: 2.34271e+07 muA
** NormalTransistorNmos: 2.34271e+07 muA
** NormalTransistorNmos: 6.74082e+08 muA
** DiodeTransistorNmos: 6.74083e+08 muA
** NormalTransistorPmos: -6.74081e+08 muA
** NormalTransistorPmos: -6.74082e+08 muA
** DiodeTransistorNmos: 2.31524e+08 muA
** NormalTransistorNmos: 2.31524e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.00499e+07 muA
** DiodeTransistorPmos: -7.56427e+08 muA


** Expected Voltages: 
** ibias: 1.29201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.08501  V
** out: 2.5  V
** outFirstStage: 4.10601  V
** outInputVoltageBiasXXnXX1: 1.32601  V
** outSourceVoltageBiasXXnXX1: 0.663001  V
** outSourceVoltageBiasXXnXX2: 0.647001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.27301  V
** out1: 3.54201  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.65001  V
** inner: 0.663001  V
** inner: 0.643001  V


.END