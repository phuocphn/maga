** Name: two_stage_single_output_op_amp_121_8

.MACRO two_stage_single_output_op_amp_121_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=7e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=5e-6
mMainBias3 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=42e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=11e-6
mTelescopicFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=78e-6
mTelescopicFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=31e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=31e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=31e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mSecondStage1StageBias11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=211e-6
mTelescopicFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=31e-6
mMainBias13 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=60e-6
mTelescopicFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=126e-6
mTelescopicFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=126e-6
mTelescopicFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=216e-6
mMainBias19 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=102e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=362e-6
mTelescopicFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=216e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.5e-12
.EOM two_stage_single_output_op_amp_121_8

** Expected Performance Values: 
** Gain: 148 dB
** Power consumption: 3.63101 mW
** Area: 7867 (mu_m)^2
** Transit frequency: 5.92201 MHz
** Transit frequency with error factor: 5.92187 MHz
** Slew rate: 7.36378 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.69001 V
** VoutMin: 0.820001 V
** VcmMax: 4.93001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 7.84801e+06 muA
** NormalTransistorNmos: 3.00231e+07 muA
** NormalTransistorPmos: -1.88589e+07 muA
** NormalTransistorNmos: 2.95221e+07 muA
** NormalTransistorNmos: 2.95221e+07 muA
** NormalTransistorPmos: -2.95229e+07 muA
** NormalTransistorPmos: -2.95239e+07 muA
** NormalTransistorPmos: -2.95229e+07 muA
** NormalTransistorPmos: -2.95239e+07 muA
** NormalTransistorNmos: 7.79011e+07 muA
** NormalTransistorNmos: 7.79001e+07 muA
** NormalTransistorNmos: 2.95221e+07 muA
** NormalTransistorNmos: 2.95221e+07 muA
** NormalTransistorNmos: 6.00478e+08 muA
** NormalTransistorNmos: 6.00477e+08 muA
** NormalTransistorPmos: -6.00477e+08 muA
** DiodeTransistorNmos: 1.88581e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.84899e+06 muA
** DiodeTransistorPmos: -3.00239e+07 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.65001  V
** out: 2.5  V
** outFirstStage: 4.13001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX0: 4.16601  V
** outVoltageBiasXXpXX1: 3.56601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.565001  V
** innerTransistorStack1Load2: 4.32501  V
** innerTransistorStack2Load2: 4.32501  V
** out1: 4.11101  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.481001  V


.END