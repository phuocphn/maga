** Name: two_stage_single_output_op_amp_76_6

.MACRO two_stage_single_output_op_amp_76_6 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=229e-6
mMainBias2 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=7e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=212e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=6e-6
mMainBias6 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=429e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=229e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=77e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=77e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=212e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mSecondStage1Transconductor15 out inputVoltageBiasXXnXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad16 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=115e-6
mMainBias17 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mMainBias18 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=70e-6
mFoldedCascodeFirstStageLoad19 FirstStageYout1 outInputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=541e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
mMainBias22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mMainBias23 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mSecondStage1StageBias24 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=429e-6
mFoldedCascodeFirstStageLoad25 outFirstStage outInputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=541e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.5e-12
.EOM two_stage_single_output_op_amp_76_6

** Expected Performance Values: 
** Gain: 179 dB
** Power consumption: 14.9811 mW
** Area: 6386 (mu_m)^2
** Transit frequency: 15.9471 MHz
** Transit frequency with error factor: 15.947 MHz
** Slew rate: 11.1789 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 3.02001 V
** VoutMin: 0.390001 V
** VcmMax: 4.66001 V
** VcmMin: 1.33001 V


** Expected Currents: 
** NormalTransistorNmos: 2.66801e+07 muA
** NormalTransistorNmos: 1.00222e+08 muA
** NormalTransistorPmos: -2.1322e+08 muA
** NormalTransistorPmos: -2.19718e+08 muA
** NormalTransistorPmos: -3.68478e+08 muA
** NormalTransistorPmos: -2.19718e+08 muA
** NormalTransistorPmos: -3.68478e+08 muA
** DiodeTransistorNmos: 2.19719e+08 muA
** NormalTransistorNmos: 2.19719e+08 muA
** NormalTransistorNmos: 2.19719e+08 muA
** NormalTransistorNmos: 2.97519e+08 muA
** DiodeTransistorNmos: 2.9752e+08 muA
** NormalTransistorNmos: 1.4876e+08 muA
** NormalTransistorNmos: 1.4876e+08 muA
** NormalTransistorNmos: 1.90908e+09 muA
** NormalTransistorNmos: 1.90908e+09 muA
** NormalTransistorPmos: -1.90907e+09 muA
** DiodeTransistorPmos: -1.90907e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 2.13221e+08 muA
** DiodeTransistorPmos: -2.66809e+07 muA
** NormalTransistorPmos: -2.66819e+07 muA
** DiodeTransistorPmos: -1.00221e+08 muA
** DiodeTransistorPmos: -1.00222e+08 muA


** Expected Voltages: 
** ibias: 1.17501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.905001  V
** out: 2.5  V
** outFirstStage: 0.598001  V
** outInputVoltageBiasXXpXX1: 2.45401  V
** outInputVoltageBiasXXpXX2: 2.37201  V
** outSourceVoltageBiasXXnXX1: 0.588001  V
** outSourceVoltageBiasXXpXX1: 3.72701  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.94401  V
** innerTransconductance: 0.306001  V
** inner: 0.586001  V
** inner: 3.72001  V


.END