** Name: two_stage_single_output_op_amp_82_5

.MACRO two_stage_single_output_op_amp_82_5 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=10e-6 W=187e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=10e-6 W=187e-6
mMainBias3 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=13e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=67e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=25e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=72e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=319e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=157e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=10e-6 W=187e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=16e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=67e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mMainBias14 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=326e-6
mSecondStage1Transconductor15 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=305e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=187e-6
mMainBias17 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=387e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=42e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=72e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=319e-6
mFoldedCascodeFirstStageLoad23 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=42e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_82_5

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 9.76401 mW
** Area: 14469 (mu_m)^2
** Transit frequency: 9.09501 MHz
** Transit frequency with error factor: 9.09503 MHz
** Slew rate: 7.76917 V/mu_s
** Phase margin: 65.3172°
** CMRR: 142 dB
** VoutMax: 3.09001 V
** VoutMin: 0.5 V
** VcmMax: 5.11001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 2.92729e+08 muA
** NormalTransistorNmos: 2.49977e+08 muA
** NormalTransistorPmos: -3.56179e+07 muA
** NormalTransistorPmos: -6.09579e+07 muA
** NormalTransistorPmos: -3.56179e+07 muA
** NormalTransistorPmos: -6.09579e+07 muA
** DiodeTransistorNmos: 3.56171e+07 muA
** NormalTransistorNmos: 3.56171e+07 muA
** NormalTransistorNmos: 3.56171e+07 muA
** DiodeTransistorNmos: 3.56171e+07 muA
** NormalTransistorNmos: 5.06781e+07 muA
** DiodeTransistorNmos: 5.06791e+07 muA
** NormalTransistorNmos: 2.53391e+07 muA
** NormalTransistorNmos: 2.53391e+07 muA
** NormalTransistorNmos: 1.27814e+09 muA
** NormalTransistorPmos: -1.27813e+09 muA
** DiodeTransistorPmos: -1.27813e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.92728e+08 muA
** NormalTransistorPmos: -2.92729e+08 muA
** DiodeTransistorPmos: -2.49976e+08 muA
** DiodeTransistorPmos: -2.49977e+08 muA


** Expected Voltages: 
** ibias: 1.18901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.82501  V
** out: 2.5  V
** outFirstStage: 0.905001  V
** outInputVoltageBiasXXpXX1: 2.52801  V
** outSourceVoltageBiasXXnXX1: 0.595001  V
** outSourceVoltageBiasXXpXX1: 3.76401  V
** outSourceVoltageBiasXXpXX2: 4.13901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 3.60601  V
** sourceGCC2: 3.60601  V
** sourceTransconductance: 1.90101  V
** inner: 0.593001  V
** inner: 3.76401  V


.END