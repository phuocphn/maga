** Name: two_stage_single_output_op_amp_21_4

.MACRO two_stage_single_output_op_amp_21_4 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=39e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=10e-6 W=76e-6
mSecondStage1StageBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=62e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=19e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=39e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=152e-6
mSecondStage1Transconductor8 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=9e-6 W=570e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=10e-6 W=76e-6
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=76e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=29e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=567e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=580e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=76e-6
mMainBias16 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=279e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_21_4

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 4.54101 mW
** Area: 11326 (mu_m)^2
** Transit frequency: 3.35201 MHz
** Transit frequency with error factor: 3.34895 MHz
** Slew rate: 6.68511 V/mu_s
** Phase margin: 69.328°
** CMRR: 100 dB
** negPSRR: 95 dB
** posPSRR: 99 dB
** VoutMax: 3.96001 V
** VoutMin: 0.690001 V
** VcmMax: 3.08001 V
** VcmMin: 0.610001 V


** Expected Currents: 
** NormalTransistorPmos: -2.82871e+08 muA
** DiodeTransistorNmos: 1.52081e+07 muA
** DiodeTransistorNmos: 1.52071e+07 muA
** NormalTransistorNmos: 1.52081e+07 muA
** NormalTransistorNmos: 1.52071e+07 muA
** NormalTransistorPmos: -3.04169e+07 muA
** NormalTransistorPmos: -3.04159e+07 muA
** NormalTransistorPmos: -1.52089e+07 muA
** NormalTransistorPmos: -1.52089e+07 muA
** NormalTransistorNmos: 5.7487e+08 muA
** NormalTransistorNmos: 5.74869e+08 muA
** NormalTransistorPmos: -5.74869e+08 muA
** NormalTransistorPmos: -5.74868e+08 muA
** DiodeTransistorNmos: 2.82872e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.46301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.772001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.09801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.619001  V
** innerStageBias: 4.26901  V
** innerTransistorStack2Load1: 0.618001  V
** out1: 1.17701  V
** sourceTransconductance: 3.38001  V
** innerStageBias: 4.26201  V
** innerTransconductance: 0.367001  V


.END