** Name: two_stage_single_output_op_amp_93_9

.MACRO two_stage_single_output_op_amp_93_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=19e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=27e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=553e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=121e-6
mTelescopicFirstStageLoad5 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=10e-6 W=16e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=22e-6
mTelescopicFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=22e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=11e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=11e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=27e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=553e-6
mTelescopicFirstStageLoad12 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=22e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=43e-6
mTelescopicFirstStageStageBias14 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=8e-6 W=319e-6
mTelescopicFirstStageLoad15 FirstStageYout1 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=10e-6 W=16e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=365e-6
mTelescopicFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=30e-6
mMainBias18 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=25e-6
mMainBias19 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=147e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.60001e-12
.EOM two_stage_single_output_op_amp_93_9

** Expected Performance Values: 
** Gain: 140 dB
** Power consumption: 3.75501 mW
** Area: 10770 (mu_m)^2
** Transit frequency: 2.63901 MHz
** Transit frequency with error factor: 2.6391 MHz
** Slew rate: 20.4087 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** VoutMax: 4.30001 V
** VoutMin: 0.700001 V
** VcmMax: 4 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorNmos: 2.23941e+07 muA
** NormalTransistorPmos: -2.59199e+07 muA
** NormalTransistorPmos: -1.52119e+08 muA
** NormalTransistorNmos: 6.98501e+06 muA
** NormalTransistorNmos: 6.98401e+06 muA
** NormalTransistorPmos: -6.98599e+06 muA
** NormalTransistorPmos: -6.98499e+06 muA
** DiodeTransistorPmos: -6.98599e+06 muA
** NormalTransistorNmos: 1.66087e+08 muA
** NormalTransistorNmos: 6.98401e+06 muA
** NormalTransistorNmos: 6.98401e+06 muA
** NormalTransistorNmos: 5.2663e+08 muA
** DiodeTransistorNmos: 5.2663e+08 muA
** NormalTransistorPmos: -5.26629e+08 muA
** DiodeTransistorNmos: 2.59191e+07 muA
** NormalTransistorNmos: 2.59181e+07 muA
** DiodeTransistorNmos: 1.5212e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.23949e+07 muA


** Expected Voltages: 
** ibias: 0.627001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.73701  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 3.71701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 3.94001  V
** out1: 3.17801  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.554001  V


.END