** Name: two_stage_single_output_op_amp_204_11

.MACRO two_stage_single_output_op_amp_204_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=51e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=51e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=9e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=104e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=36e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=6e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=11e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=51e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=14e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=36e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=512e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=104e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=528e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=7e-6 W=51e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=14e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=15e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mSimpleFirstStageLoad19 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=354e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=584e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=578e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=354e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=120e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.40001e-12
.EOM two_stage_single_output_op_amp_204_11

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 5.28701 mW
** Area: 14984 (mu_m)^2
** Transit frequency: 4.34701 MHz
** Transit frequency with error factor: 4.32028 MHz
** Slew rate: 4.0965 V/mu_s
** Phase margin: 60.1606°
** CMRR: 95 dB
** VoutMax: 4.34001 V
** VoutMin: 0.710001 V
** VcmMax: 4.87001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 1.50111e+07 muA
** NormalTransistorNmos: 7.00501e+06 muA
** NormalTransistorPmos: -7.69189e+07 muA
** DiodeTransistorNmos: 2.09446e+08 muA
** NormalTransistorNmos: 2.09447e+08 muA
** NormalTransistorNmos: 2.09446e+08 muA
** DiodeTransistorNmos: 2.09447e+08 muA
** NormalTransistorPmos: -2.22778e+08 muA
** NormalTransistorPmos: -2.22778e+08 muA
** NormalTransistorNmos: 2.66651e+07 muA
** DiodeTransistorNmos: 2.66641e+07 muA
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 5.02823e+08 muA
** NormalTransistorNmos: 5.02822e+08 muA
** NormalTransistorPmos: -5.02822e+08 muA
** NormalTransistorPmos: -5.02823e+08 muA
** DiodeTransistorNmos: 7.69181e+07 muA
** NormalTransistorNmos: 7.69171e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.50119e+07 muA
** DiodeTransistorPmos: -7.00599e+06 muA


** Expected Voltages: 
** ibias: 1.125  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.21601  V
** outInputVoltageBiasXXnXX1: 1.22801  V
** outSourceVoltageBiasXXnXX1: 0.614001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 3.90301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.10501  V
** innerTransistorStack1Load1: 1.10501  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.570001  V
** innerTransconductance: 4.69001  V
** inner: 0.613001  V


.END