** Name: two_stage_single_output_op_amp_151_7

.MACRO two_stage_single_output_op_amp_151_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=5e-6 W=8e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=23e-6
mSimpleFirstStageTransconductor5 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=101e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=73e-6
mMainBias8 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=32e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=8e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=101e-6
mSimpleFirstStageLoad12 FirstStageYinnerOutputLoad1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=109e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=361e-6
mSimpleFirstStageLoad14 outFirstStage inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=109e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.2001e-12
.EOM two_stage_single_output_op_amp_151_7

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 3.14901 mW
** Area: 5743 (mu_m)^2
** Transit frequency: 4.16401 MHz
** Transit frequency with error factor: 4.1523 MHz
** Slew rate: 3.92454 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.75 V
** VoutMin: 0.150001 V
** VcmMax: 4.85001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorNmos: 2.13121e+07 muA
** DiodeTransistorNmos: 7.50291e+07 muA
** NormalTransistorNmos: 7.50281e+07 muA
** NormalTransistorNmos: 7.50291e+07 muA
** DiodeTransistorNmos: 7.50281e+07 muA
** NormalTransistorPmos: -9.90759e+07 muA
** NormalTransistorPmos: -9.90759e+07 muA
** NormalTransistorNmos: 4.80911e+07 muA
** NormalTransistorNmos: 2.40461e+07 muA
** NormalTransistorNmos: 2.40461e+07 muA
** NormalTransistorNmos: 4.00318e+08 muA
** NormalTransistorPmos: -4.00317e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.13129e+07 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.88101  V
** out: 2.5  V
** outFirstStage: 4.18601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.30501  V
** innerSourceLoad1: 1.15201  V
** innerTransistorStack1Load1: 1.15201  V
** sourceTransconductance: 1.94501  V


.END