** Name: two_stage_single_output_op_amp_80_7

.MACRO two_stage_single_output_op_amp_80_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mMainBias2 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=29e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=5e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=81e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=20e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=25e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=51e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=68e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=68e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=81e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=1e-6 W=284e-6
mFoldedCascodeFirstStageLoad15 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=51e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=283e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=143e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=143e-6
mMainBias19 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=195e-6
mMainBias20 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=405e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=319e-6
mFoldedCascodeFirstStageLoad22 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=283e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=6e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.60001e-12
.EOM two_stage_single_output_op_amp_80_7

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 10.0011 mW
** Area: 8044 (mu_m)^2
** Transit frequency: 4.65901 MHz
** Transit frequency with error factor: 4.65902 MHz
** Slew rate: 4.97685 V/mu_s
** Phase margin: 60.1606°
** CMRR: 147 dB
** VoutMax: 4.25 V
** VoutMin: 0.260001 V
** VcmMax: 5.15001 V
** VcmMin: 1.33001 V


** Expected Currents: 
** NormalTransistorPmos: -2.43999e+06 muA
** NormalTransistorPmos: -7.88429e+07 muA
** NormalTransistorPmos: -1.63044e+08 muA
** NormalTransistorPmos: -3.83119e+07 muA
** NormalTransistorPmos: -5.81629e+07 muA
** NormalTransistorPmos: -3.83119e+07 muA
** NormalTransistorPmos: -5.81629e+07 muA
** NormalTransistorNmos: 3.83111e+07 muA
** NormalTransistorNmos: 3.83101e+07 muA
** NormalTransistorNmos: 3.83111e+07 muA
** NormalTransistorNmos: 3.83101e+07 muA
** NormalTransistorNmos: 3.96991e+07 muA
** DiodeTransistorNmos: 3.96981e+07 muA
** NormalTransistorNmos: 1.98501e+07 muA
** NormalTransistorNmos: 1.98501e+07 muA
** NormalTransistorNmos: 1.61947e+09 muA
** NormalTransistorPmos: -1.61946e+09 muA
** DiodeTransistorNmos: 2.43901e+06 muA
** NormalTransistorNmos: 2.43801e+06 muA
** DiodeTransistorNmos: 7.88421e+07 muA
** DiodeTransistorNmos: 1.63045e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.943001  V
** inputVoltageBiasXXnXX3: 0.664001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.15001  V
** outSourceVoltageBiasXXnXX1: 0.575001  V
** outSourceVoltageBiasXXpXX1: 4.17601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.91801  V
** inner: 0.575001  V


.END