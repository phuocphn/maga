** Name: symmetrical_op_amp196

.MACRO symmetrical_op_amp196 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=9e-6
mSecondStage1StageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=44e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=1e-6 W=44e-6
mSymmetricalFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=247e-6
mMainBias5 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=247e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias7 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=44e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=62e-6
mSecondStage1StageBias10 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=1e-6 W=44e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=62e-6
mMainBias12 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=89e-6
mSymmetricalFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=42e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=42e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=40e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=40e-6
mSymmetricalFirstStageLoad17 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=335e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=317e-6
mSecondStage1Transconductor19 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=317e-6
mSymmetricalFirstStageLoad20 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=335e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp196

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 3.19401 mW
** Area: 3144 (mu_m)^2
** Transit frequency: 12.7481 MHz
** Transit frequency with error factor: 12.7478 MHz
** Slew rate: 12.8244 V/mu_s
** Phase margin: 83.6519°
** CMRR: 143 dB
** negPSRR: 128 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 0.770001 V
** VcmMax: 4.81001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 9.97591e+07 muA
** NormalTransistorPmos: -1.35822e+08 muA
** NormalTransistorPmos: -1.35823e+08 muA
** NormalTransistorPmos: -1.35822e+08 muA
** NormalTransistorPmos: -1.35823e+08 muA
** NormalTransistorNmos: 2.71646e+08 muA
** DiodeTransistorNmos: 2.71647e+08 muA
** NormalTransistorNmos: 1.35823e+08 muA
** NormalTransistorNmos: 1.35823e+08 muA
** NormalTransistorNmos: 1.28745e+08 muA
** DiodeTransistorNmos: 1.28744e+08 muA
** NormalTransistorPmos: -1.28744e+08 muA
** NormalTransistorPmos: -1.28745e+08 muA
** DiodeTransistorNmos: 1.28745e+08 muA
** NormalTransistorNmos: 1.28744e+08 muA
** NormalTransistorPmos: -1.28744e+08 muA
** NormalTransistorPmos: -1.28745e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.97599e+07 muA


** Expected Voltages: 
** ibias: 1.13301  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 0.590001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 1.18001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.567001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.93401  V
** innerTransconductance: 4.40001  V
** inner: 0.589001  V
** inner: 4.40001  V
** inner: 0.566001  V


.END