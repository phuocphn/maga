** Name: two_stage_single_output_op_amp_77_3

.MACRO two_stage_single_output_op_amp_77_3 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=48e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=49e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=42e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=8e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=88e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=49e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=31e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=31e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=75e-6
mMainBias12 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=213e-6
mSecondStage1Transconductor13 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=147e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=48e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerOutputLoad2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=83e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=162e-6
mSecondStage1StageBias19 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=340e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=83e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_77_3

** Expected Performance Values: 
** Gain: 132 dB
** Power consumption: 4.55901 mW
** Area: 8274 (mu_m)^2
** Transit frequency: 3.94601 MHz
** Transit frequency with error factor: 3.94568 MHz
** Slew rate: 3.71526 V/mu_s
** Phase margin: 69.328°
** CMRR: 149 dB
** VoutMax: 3.17001 V
** VoutMin: 0.510001 V
** VcmMax: 4.66001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 4.06121e+07 muA
** NormalTransistorPmos: -1.68539e+07 muA
** NormalTransistorPmos: -2.52899e+07 muA
** NormalTransistorPmos: -1.68539e+07 muA
** NormalTransistorPmos: -2.52899e+07 muA
** DiodeTransistorNmos: 1.68531e+07 muA
** DiodeTransistorNmos: 1.68521e+07 muA
** NormalTransistorNmos: 1.68531e+07 muA
** NormalTransistorNmos: 1.68521e+07 muA
** NormalTransistorNmos: 1.68691e+07 muA
** NormalTransistorNmos: 1.68681e+07 muA
** NormalTransistorNmos: 8.43501e+06 muA
** NormalTransistorNmos: 8.43501e+06 muA
** NormalTransistorNmos: 8.10585e+08 muA
** NormalTransistorPmos: -8.10584e+08 muA
** NormalTransistorPmos: -8.10585e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -4.06129e+07 muA
** DiodeTransistorPmos: -4.06129e+07 muA


** Expected Voltages: 
** ibias: 1.12701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.918001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.12301  V
** innerStageBias: 0.559001  V
** innerTransistorStack1Load2: 0.561001  V
** innerTransistorStack2Load2: 0.560001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 3.45001  V


.END