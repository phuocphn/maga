** Name: two_stage_single_output_op_amp_86_3

.MACRO two_stage_single_output_op_amp_86_3 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=28e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=98e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=72e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=28e-6
mMainBias7 inputVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=447e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=442e-6
mTelescopicFirstStageLoad9 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=28e-6
mMainBias10 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=105e-6
mTelescopicFirstStageLoad11 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=10e-6 W=11e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=27e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=27e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=470e-6
mMainBias15 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=61e-6
mSecondStage1StageBias16 out inputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=595e-6
mTelescopicFirstStageLoad17 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=10e-6 W=11e-6
mTelescopicFirstStageStageBias18 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=77e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_86_3

** Expected Performance Values: 
** Gain: 142 dB
** Power consumption: 4.59501 mW
** Area: 10584 (mu_m)^2
** Transit frequency: 2.55301 MHz
** Transit frequency with error factor: 2.55284 MHz
** Slew rate: 16.6387 V/mu_s
** Phase margin: 60.1606°
** CMRR: 130 dB
** VoutMax: 4.37001 V
** VoutMin: 0.300001 V
** VcmMax: 3.94001 V
** VcmMin: 0.690001 V


** Expected Currents: 
** NormalTransistorNmos: 6.66001e+07 muA
** NormalTransistorNmos: 2.82039e+08 muA
** NormalTransistorPmos: -6.21529e+07 muA
** NormalTransistorPmos: -5.92699e+06 muA
** NormalTransistorPmos: -5.92699e+06 muA
** NormalTransistorNmos: 5.92601e+06 muA
** NormalTransistorNmos: 5.92601e+06 muA
** DiodeTransistorNmos: 5.92601e+06 muA
** NormalTransistorPmos: -7.84559e+07 muA
** NormalTransistorPmos: -5.92799e+06 muA
** NormalTransistorPmos: -5.92799e+06 muA
** NormalTransistorNmos: 4.76292e+08 muA
** NormalTransistorPmos: -4.76291e+08 muA
** NormalTransistorPmos: -4.76292e+08 muA
** DiodeTransistorNmos: 6.21521e+07 muA
** DiodeTransistorPmos: -6.66009e+07 muA
** DiodeTransistorPmos: -2.82038e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.10001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.598001  V
** inputVoltageBiasXXpXX2: 1.93601  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outVoltageBiasXXpXX1: 1.93301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.22001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 3.04401  V
** sourceGCC2: 3.04401  V
** innerStageBias: 2.79801  V


.END