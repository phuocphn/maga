** Name: two_stage_single_output_op_amp_147_9

.MACRO two_stage_single_output_op_amp_147_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=11e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=7e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=456e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=46e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=30e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=456e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=11e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=30e-6
mSimpleFirstStageLoad14 FirstStageYinnerOutputLoad1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=419e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=101e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=144e-6
mSimpleFirstStageLoad17 outFirstStage ibias sourcePmos sourcePmos pmos4 L=3e-6 W=419e-6
mMainBias18 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=240e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.5e-12
.EOM two_stage_single_output_op_amp_147_9

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 8.69601 mW
** Area: 9750 (mu_m)^2
** Transit frequency: 4.15001 MHz
** Transit frequency with error factor: 4.14135 MHz
** Slew rate: 3.91108 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 1.35001 V
** VcmMax: 5.21001 V
** VcmMin: 0.770001 V


** Expected Currents: 
** NormalTransistorPmos: -2.21689e+07 muA
** NormalTransistorPmos: -5.26799e+07 muA
** DiodeTransistorNmos: 6.25241e+07 muA
** DiodeTransistorNmos: 6.25251e+07 muA
** NormalTransistorNmos: 6.25241e+07 muA
** NormalTransistorNmos: 6.25251e+07 muA
** NormalTransistorPmos: -9.10949e+07 muA
** NormalTransistorPmos: -9.10949e+07 muA
** NormalTransistorNmos: 5.71391e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 1.46209e+09 muA
** DiodeTransistorNmos: 1.46209e+09 muA
** NormalTransistorPmos: -1.46208e+09 muA
** DiodeTransistorNmos: 2.21681e+07 muA
** NormalTransistorNmos: 2.21671e+07 muA
** DiodeTransistorNmos: 5.26791e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.76001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.880001  V
** outVoltageBiasXXnXX2: 0.624001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.19501  V
** innerSourceLoad1: 1.15301  V
** innerTransistorStack2Load1: 1.15301  V
** sourceTransconductance: 1.94501  V
** inner: 0.879001  V


.END