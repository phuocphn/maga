** Name: two_stage_single_output_op_amp_79_12

.MACRO two_stage_single_output_op_amp_79_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=151e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=49e-6
mMainBias3 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=165e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=444e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=40e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=42e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=113e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=113e-6
mFoldedCascodeFirstStageLoad10 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=96e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=17e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=180e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=151e-6
mSecondStage1StageBias15 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=444e-6
mFoldedCascodeFirstStageLoad16 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=96e-6
mMainBias17 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=132e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=176e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=127e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=127e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mMainBias22 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=513e-6
mMainBias23 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=309e-6
mMainBias24 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=373e-6
mSecondStage1Transconductor25 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=582e-6
mFoldedCascodeFirstStageLoad26 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=176e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.9001e-12
.EOM two_stage_single_output_op_amp_79_12

** Expected Performance Values: 
** Gain: 175 dB
** Power consumption: 11.1311 mW
** Area: 10534 (mu_m)^2
** Transit frequency: 4.58901 MHz
** Transit frequency with error factor: 4.58882 MHz
** Slew rate: 3.59968 V/mu_s
** Phase margin: 64.7443°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 0.870001 V
** VcmMax: 5.21001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 2.03068e+08 muA
** NormalTransistorPmos: -3.48504e+08 muA
** NormalTransistorPmos: -2.06299e+08 muA
** NormalTransistorPmos: -2.49613e+08 muA
** NormalTransistorPmos: -5.38989e+07 muA
** NormalTransistorPmos: -8.62769e+07 muA
** NormalTransistorPmos: -5.38989e+07 muA
** NormalTransistorPmos: -8.62769e+07 muA
** NormalTransistorNmos: 5.38981e+07 muA
** NormalTransistorNmos: 5.38971e+07 muA
** NormalTransistorNmos: 5.38981e+07 muA
** NormalTransistorNmos: 5.38971e+07 muA
** NormalTransistorNmos: 6.47571e+07 muA
** NormalTransistorNmos: 6.47561e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 1.02619e+09 muA
** DiodeTransistorNmos: 1.02619e+09 muA
** NormalTransistorPmos: -1.02618e+09 muA
** NormalTransistorPmos: -1.02618e+09 muA
** DiodeTransistorNmos: 3.48505e+08 muA
** NormalTransistorNmos: 3.48504e+08 muA
** DiodeTransistorNmos: 2.063e+08 muA
** DiodeTransistorNmos: 2.49614e+08 muA
** DiodeTransistorPmos: -2.03067e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.27601  V
** inputVoltageBiasXXnXX2: 0.954001  V
** inputVoltageBiasXXnXX3: 0.595001  V
** out: 2.5  V
** outFirstStage: 4.12801  V
** outSourceVoltageBiasXXnXX1: 0.638001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.390001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.43501  V
** sourceGCC2: 4.43501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.69201  V
** inner: 0.637001  V


.END