** Name: two_stage_single_output_op_amp_61_1

.MACRO two_stage_single_output_op_amp_61_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=7e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=11e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=16e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=95e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=95e-6
mMainBias9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=29e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=74e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=16e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=48e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=119e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=119e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=8e-6 W=210e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=523e-6
mFoldedCascodeFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=8e-6 W=231e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.5e-12
.EOM two_stage_single_output_op_amp_61_1

** Expected Performance Values: 
** Gain: 118 dB
** Power consumption: 3.56201 mW
** Area: 7106 (mu_m)^2
** Transit frequency: 3.39901 MHz
** Transit frequency with error factor: 3.39892 MHz
** Slew rate: 3.97218 V/mu_s
** Phase margin: 60.1606°
** CMRR: 141 dB
** VoutMax: 4.75 V
** VoutMin: 0.610001 V
** VcmMax: 3.18001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.38091e+07 muA
** NormalTransistorNmos: 2.30861e+07 muA
** NormalTransistorNmos: 2.99721e+07 muA
** NormalTransistorNmos: 4.52351e+07 muA
** NormalTransistorNmos: 2.99721e+07 muA
** NormalTransistorNmos: 4.52351e+07 muA
** DiodeTransistorPmos: -2.99729e+07 muA
** NormalTransistorPmos: -2.99729e+07 muA
** NormalTransistorPmos: -2.99729e+07 muA
** NormalTransistorPmos: -3.05289e+07 muA
** NormalTransistorPmos: -3.05299e+07 muA
** NormalTransistorPmos: -1.52639e+07 muA
** NormalTransistorPmos: -1.52639e+07 muA
** NormalTransistorNmos: 5.7506e+08 muA
** NormalTransistorPmos: -5.75059e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.38099e+07 muA
** DiodeTransistorPmos: -2.30869e+07 muA


** Expected Voltages: 
** ibias: 1.21901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 1.01401  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX2: 4.18801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.50401  V
** innerTransistorStack2Load2: 4.49001  V
** out1: 4.27101  V
** sourceGCC1: 0.515001  V
** sourceGCC2: 0.515001  V
** sourceTransconductance: 3.25301  V


.END