** Name: two_stage_single_output_op_amp_32_10

.MACRO two_stage_single_output_op_amp_32_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=14e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=41e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=501e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=165e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=41e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mMainBias10 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=579e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=165e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=51e-6
mSimpleFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=501e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=353e-6
mSecondStage1Transconductor16 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=7e-6 W=359e-6
mMainBias18 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=28e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18e-12
.EOM two_stage_single_output_op_amp_32_10

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 7.02601 mW
** Area: 14976 (mu_m)^2
** Transit frequency: 6.12201 MHz
** Transit frequency with error factor: 6.11891 MHz
** Slew rate: 5.76978 V/mu_s
** Phase margin: 60.1606°
** CMRR: 106 dB
** negPSRR: 110 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 0.310001 V
** VcmMax: 4.42001 V
** VcmMin: 1.81001 V


** Expected Currents: 
** NormalTransistorNmos: 9.88801e+06 muA
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -3.51589e+07 muA
** NormalTransistorPmos: -5.23789e+07 muA
** NormalTransistorPmos: -5.23789e+07 muA
** DiodeTransistorPmos: -5.23789e+07 muA
** NormalTransistorNmos: 1.04756e+08 muA
** DiodeTransistorNmos: 1.04755e+08 muA
** NormalTransistorNmos: 5.23781e+07 muA
** NormalTransistorNmos: 5.23781e+07 muA
** NormalTransistorNmos: 1.14395e+09 muA
** NormalTransistorPmos: -1.14394e+09 muA
** NormalTransistorPmos: -1.14395e+09 muA
** DiodeTransistorNmos: 3.51581e+07 muA
** NormalTransistorNmos: 3.51581e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.88899e+06 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 0.711001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.68901  V
** out: 2.5  V
** outFirstStage: 4.01101  V
** outInputVoltageBiasXXnXX1: 1.65801  V
** outSourceVoltageBiasXXnXX1: 0.829001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.24901  V
** out1: 3.44701  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.57501  V
** inner: 0.829001  V


.END