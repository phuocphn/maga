** Name: one_stage_single_output_op_amp90

.MACRO one_stage_single_output_op_amp90 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=23e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=29e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=6e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mTelescopicFirstStageLoad7 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=23e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=6e-6 W=208e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=222e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=222e-6
mTelescopicFirstStageLoad12 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=6e-6 W=208e-6
mMainBias13 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=14e-6
mTelescopicFirstStageStageBias14 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=268e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp90

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 0.595001 mW
** Area: 4783 (mu_m)^2
** Transit frequency: 4.74301 MHz
** Transit frequency with error factor: 4.74345 MHz
** Slew rate: 4.6913 V/mu_s
** Phase margin: 64.7443°
** CMRR: 151 dB
** VoutMax: 4.30001 V
** VoutMin: 0.710001 V
** VcmMax: 4.01001 V
** VcmMin: 0.820001 V


** Expected Currents: 
** NormalTransistorNmos: 3.97701e+06 muA
** NormalTransistorPmos: -4.91699e+06 muA
** NormalTransistorPmos: -4.50799e+07 muA
** NormalTransistorPmos: -4.50819e+07 muA
** DiodeTransistorNmos: 4.50791e+07 muA
** NormalTransistorNmos: 4.50801e+07 muA
** NormalTransistorNmos: 4.50811e+07 muA
** DiodeTransistorNmos: 4.50801e+07 muA
** NormalTransistorPmos: -9.41389e+07 muA
** NormalTransistorPmos: -4.50809e+07 muA
** NormalTransistorPmos: -4.50809e+07 muA
** DiodeTransistorNmos: 4.91601e+06 muA
** DiodeTransistorPmos: -3.97799e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.15701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outVoltageBiasXXnXX0: 0.592001  V
** outVoltageBiasXXpXX1: 2.18001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21401  V
** innerTransistorStack1Load2: 0.557001  V
** innerTransistorStack2Load2: 0.557001  V
** out1: 1.11401  V
** sourceGCC1: 3.01501  V
** sourceGCC2: 3.01501  V


.END