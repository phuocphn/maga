** Name: two_stage_single_output_op_amp_143_11

.MACRO two_stage_single_output_op_amp_143_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=118e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mSecondStage1StageBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=90e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=185e-6
mSimpleFirstStageLoad7 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=118e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=49e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=598e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=240e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=14e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=185e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=49e-6
mMainBias14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=80e-6
mSimpleFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=243e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=567e-6
mMainBias17 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=61e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad19 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=243e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.7001e-12
.EOM two_stage_single_output_op_amp_143_11

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 14.9271 mW
** Area: 10423 (mu_m)^2
** Transit frequency: 10.6711 MHz
** Transit frequency with error factor: 10.608 MHz
** Slew rate: 10.1691 V/mu_s
** Phase margin: 60.1606°
** CMRR: 94 dB
** VoutMax: 4.25 V
** VoutMin: 0.720001 V
** VcmMax: 4.91001 V
** VcmMin: 0.900001 V


** Expected Currents: 
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorNmos: 1.96061e+08 muA
** NormalTransistorPmos: -1.33347e+08 muA
** NormalTransistorNmos: 4.68671e+08 muA
** NormalTransistorNmos: 4.68672e+08 muA
** DiodeTransistorNmos: 4.68671e+08 muA
** NormalTransistorPmos: -5.28713e+08 muA
** NormalTransistorPmos: -5.28713e+08 muA
** NormalTransistorNmos: 1.20088e+08 muA
** NormalTransistorNmos: 6.00431e+07 muA
** NormalTransistorNmos: 6.00431e+07 muA
** NormalTransistorNmos: 1.46669e+09 muA
** NormalTransistorNmos: 1.46669e+09 muA
** NormalTransistorPmos: -1.46668e+09 muA
** NormalTransistorPmos: -1.46668e+09 muA
** DiodeTransistorNmos: 1.33348e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.21839e+08 muA
** DiodeTransistorPmos: -1.9606e+08 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.12601  V
** out: 2.5  V
** outFirstStage: 4.05401  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 3.94101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 1.05801  V
** out1: 2.09501  V
** sourceTransconductance: 1.94301  V
** innerStageBias: 0.342001  V
** innerTransconductance: 4.61801  V


.END