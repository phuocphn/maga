** Name: two_stage_single_output_op_amp_75_5

.MACRO two_stage_single_output_op_amp_75_5 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=71e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=4e-6 W=4e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=4e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=499e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=71e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=60e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=60e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=127e-6
mMainBias13 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSecondStage1Transconductor14 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=482e-6
mFoldedCascodeFirstStageLoad15 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=123e-6
mMainBias16 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=421e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=28e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=28e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=499e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=421e-6
mMainBias23 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=12e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.4001e-12
.EOM two_stage_single_output_op_amp_75_5

** Expected Performance Values: 
** Gain: 142 dB
** Power consumption: 8.44901 mW
** Area: 10272 (mu_m)^2
** Transit frequency: 5.25801 MHz
** Transit frequency with error factor: 5.25805 MHz
** Slew rate: 3.67995 V/mu_s
** Phase margin: 60.1606°
** CMRR: 144 dB
** VoutMax: 3.02001 V
** VoutMin: 0.190001 V
** VcmMax: 4.66001 V
** VcmMin: 1.35001 V


** Expected Currents: 
** NormalTransistorNmos: 1.18401e+07 muA
** NormalTransistorNmos: 1.00651e+07 muA
** NormalTransistorPmos: -3.02709e+07 muA
** NormalTransistorPmos: -4.24619e+07 muA
** NormalTransistorPmos: -7.10729e+07 muA
** NormalTransistorPmos: -4.24619e+07 muA
** NormalTransistorPmos: -7.10729e+07 muA
** DiodeTransistorNmos: 4.24611e+07 muA
** NormalTransistorNmos: 4.24611e+07 muA
** NormalTransistorNmos: 4.24611e+07 muA
** NormalTransistorNmos: 5.72251e+07 muA
** NormalTransistorNmos: 5.72261e+07 muA
** NormalTransistorNmos: 2.86121e+07 muA
** NormalTransistorNmos: 2.86121e+07 muA
** NormalTransistorNmos: 1.48558e+09 muA
** NormalTransistorPmos: -1.48557e+09 muA
** DiodeTransistorPmos: -1.48557e+09 muA
** DiodeTransistorNmos: 3.02701e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.18389e+07 muA
** NormalTransistorPmos: -1.18379e+07 muA
** DiodeTransistorPmos: -1.00659e+07 muA
** DiodeTransistorPmos: -1.00669e+07 muA


** Expected Voltages: 
** ibias: 0.622001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.595001  V
** outInputVoltageBiasXXpXX1: 2.45401  V
** outSourceVoltageBiasXXpXX1: 3.72801  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX1: 1  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.417001  V
** innerTransistorStack2Load2: 0.438001  V
** out1: 0.627001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.94501  V
** inner: 3.72001  V


.END