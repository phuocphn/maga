** Name: two_stage_single_output_op_amp_105_7

.MACRO two_stage_single_output_op_amp_105_7 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=24e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=7e-6 W=17e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=8e-6 W=83e-6
mMainBias5 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=156e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=64e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=24e-6
mMainBias8 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=17e-6
mMainBias11 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=99e-6
mTelescopicFirstStageStageBias12 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=570e-6
mTelescopicFirstStageLoad13 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=16e-6
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=59e-6
mTelescopicFirstStageTransconductor15 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=59e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=122e-6
mTelescopicFirstStageLoad17 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=16e-6
mTelescopicFirstStageStageBias18 sourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=8e-6 W=570e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_105_7

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 5.32801 mW
** Area: 14496 (mu_m)^2
** Transit frequency: 2.62001 MHz
** Transit frequency with error factor: 2.61984 MHz
** Slew rate: 34.102 V/mu_s
** Phase margin: 60.1606°
** CMRR: 130 dB
** VoutMax: 3.46001 V
** VoutMin: 0.180001 V
** VcmMax: 3 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 1.40708e+08 muA
** NormalTransistorNmos: 4.28721e+07 muA
** NormalTransistorPmos: -6.53099e+06 muA
** NormalTransistorPmos: -6.53099e+06 muA
** DiodeTransistorNmos: 6.53001e+06 muA
** DiodeTransistorNmos: 6.53101e+06 muA
** NormalTransistorNmos: 6.53001e+06 muA
** NormalTransistorNmos: 6.53101e+06 muA
** NormalTransistorPmos: -1.53772e+08 muA
** NormalTransistorPmos: -1.53773e+08 muA
** NormalTransistorPmos: -6.53199e+06 muA
** NormalTransistorPmos: -6.53199e+06 muA
** NormalTransistorNmos: 8.59044e+08 muA
** NormalTransistorPmos: -8.59043e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.40707e+08 muA
** DiodeTransistorPmos: -4.28729e+07 muA
** DiodeTransistorPmos: -4.28719e+07 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.04001  V
** out: 2.5  V
** outFirstStage: 2.89101  V
** outSourceVoltageBiasXXpXX2: 4.08701  V
** outVoltageBiasXXpXX1: 2.32701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.24001  V
** innerStageBias: 3.95001  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.554001  V
** out1: 1.13801  V
** sourceGCC1: 3.04201  V
** sourceGCC2: 3.04201  V


.END