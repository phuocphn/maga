** Name: two_stage_single_output_op_amp_80_5

.MACRO two_stage_single_output_op_amp_80_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=30e-6
mFoldedCascodeFirstStageStageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=162e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=15e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=10e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=5e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=568e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=139e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=26e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=26e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=162e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
mMainBias15 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=154e-6
mSecondStage1Transconductor16 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=219e-6
mFoldedCascodeFirstStageLoad17 outFirstStage outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=139e-6
mMainBias18 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=26e-6
mFoldedCascodeFirstStageLoad19 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=245e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mMainBias22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
mSecondStage1StageBias23 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=568e-6
mFoldedCascodeFirstStageLoad24 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=245e-6
mMainBias25 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.60001e-12
.EOM two_stage_single_output_op_amp_80_5

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 6.27301 mW
** Area: 13054 (mu_m)^2
** Transit frequency: 8.12101 MHz
** Transit frequency with error factor: 8.12085 MHz
** Slew rate: 7.39323 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 3.18001 V
** VoutMin: 0.330001 V
** VcmMax: 4.66001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorNmos: 8.66501e+06 muA
** NormalTransistorNmos: 5.07661e+07 muA
** NormalTransistorPmos: -4.55459e+07 muA
** NormalTransistorPmos: -4.95659e+07 muA
** NormalTransistorPmos: -7.61499e+07 muA
** NormalTransistorPmos: -4.95659e+07 muA
** NormalTransistorPmos: -7.61499e+07 muA
** NormalTransistorNmos: 4.95651e+07 muA
** NormalTransistorNmos: 4.95641e+07 muA
** NormalTransistorNmos: 4.95651e+07 muA
** NormalTransistorNmos: 4.95641e+07 muA
** NormalTransistorNmos: 5.31711e+07 muA
** DiodeTransistorNmos: 5.31721e+07 muA
** NormalTransistorNmos: 2.65851e+07 muA
** NormalTransistorNmos: 2.65851e+07 muA
** NormalTransistorNmos: 9.87343e+08 muA
** NormalTransistorPmos: -9.87342e+08 muA
** DiodeTransistorPmos: -9.87343e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 4.55451e+07 muA
** DiodeTransistorPmos: -8.66599e+06 muA
** NormalTransistorPmos: -8.66699e+06 muA
** DiodeTransistorPmos: -5.07669e+07 muA
** DiodeTransistorPmos: -5.07669e+07 muA


** Expected Voltages: 
** ibias: 1.16301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.733001  V
** outInputVoltageBiasXXpXX1: 2.62001  V
** outSourceVoltageBiasXXnXX1: 0.582001  V
** outSourceVoltageBiasXXpXX1: 3.81001  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX2: 0.938001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.93901  V
** inner: 0.580001  V
** inner: 3.80401  V


.END