** Name: two_stage_single_output_op_amp_80_9

.MACRO two_stage_single_output_op_amp_80_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=45e-6
mMainBias2 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=8e-6
mFoldedCascodeFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=77e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=241e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=9e-6 W=24e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=33e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=27e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=107e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=48e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=48e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=42e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=42e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=77e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=45e-6
mMainBias15 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mSecondStage1StageBias16 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=241e-6
mFoldedCascodeFirstStageLoad17 outFirstStage outVoltageBiasXXnXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=107e-6
mFoldedCascodeFirstStageLoad18 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=227e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=98e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=98e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=521e-6
mFoldedCascodeFirstStageLoad22 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=227e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=44e-6
mMainBias24 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=157e-6
mMainBias25 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=149e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.40001e-12
.EOM two_stage_single_output_op_amp_80_9

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 9.94101 mW
** Area: 12203 (mu_m)^2
** Transit frequency: 3.85201 MHz
** Transit frequency with error factor: 3.85219 MHz
** Slew rate: 3.55055 V/mu_s
** Phase margin: 60.1606°
** CMRR: 147 dB
** VoutMax: 4.25 V
** VoutMin: 1.42001 V
** VcmMax: 5.12001 V
** VcmMin: 1.33001 V


** Expected Currents: 
** NormalTransistorPmos: -1.62629e+07 muA
** NormalTransistorPmos: -5.86119e+07 muA
** NormalTransistorPmos: -5.60999e+07 muA
** NormalTransistorPmos: -2.30479e+07 muA
** NormalTransistorPmos: -3.69359e+07 muA
** NormalTransistorPmos: -2.30479e+07 muA
** NormalTransistorPmos: -3.69359e+07 muA
** NormalTransistorNmos: 2.30471e+07 muA
** NormalTransistorNmos: 2.30461e+07 muA
** NormalTransistorNmos: 2.30471e+07 muA
** NormalTransistorNmos: 2.30461e+07 muA
** NormalTransistorNmos: 2.77731e+07 muA
** DiodeTransistorNmos: 2.77721e+07 muA
** NormalTransistorNmos: 1.38871e+07 muA
** NormalTransistorNmos: 1.38871e+07 muA
** NormalTransistorNmos: 1.76331e+09 muA
** DiodeTransistorNmos: 1.76331e+09 muA
** NormalTransistorPmos: -1.7633e+09 muA
** DiodeTransistorNmos: 1.62621e+07 muA
** NormalTransistorNmos: 1.62611e+07 muA
** DiodeTransistorNmos: 5.86111e+07 muA
** NormalTransistorNmos: 5.86101e+07 muA
** DiodeTransistorNmos: 5.60991e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.15401  V
** outInputVoltageBiasXXnXX2: 1.82401  V
** outSourceVoltageBiasXXnXX1: 0.577001  V
** outSourceVoltageBiasXXnXX2: 0.912001  V
** outSourceVoltageBiasXXpXX1: 4.14701  V
** outVoltageBiasXXnXX3: 0.906001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.91801  V
** inner: 0.576001  V
** inner: 0.907001  V


.END