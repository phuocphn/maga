** Name: two_stage_single_output_op_amp_38_11

.MACRO two_stage_single_output_op_amp_38_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=190e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=124e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=49e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=30e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=65e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=124e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=506e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=190e-6
mSecondStage1StageBias11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=127e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=65e-6
mMainBias13 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=22e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=61e-6
mSimpleFirstStageLoad15 FirstStageYinnerSourceLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=5e-6 W=125e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=22e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=22e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=378e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=5e-6 W=600e-6
mSimpleFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=5e-6 W=125e-6
mMainBias21 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=105e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8e-12
.EOM two_stage_single_output_op_amp_38_11

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 3.33801 mW
** Area: 14824 (mu_m)^2
** Transit frequency: 4.07701 MHz
** Transit frequency with error factor: 4.07551 MHz
** Slew rate: 3.84243 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** negPSRR: 104 dB
** posPSRR: 98 dB
** VoutMax: 4.25 V
** VoutMin: 0.860001 V
** VcmMax: 4.84001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 2.16401e+07 muA
** NormalTransistorNmos: 6.09191e+07 muA
** NormalTransistorPmos: -4.70119e+07 muA
** NormalTransistorPmos: -1.54769e+07 muA
** NormalTransistorPmos: -1.54779e+07 muA
** NormalTransistorPmos: -1.54769e+07 muA
** NormalTransistorPmos: -1.54779e+07 muA
** NormalTransistorNmos: 3.09511e+07 muA
** DiodeTransistorNmos: 3.09501e+07 muA
** NormalTransistorNmos: 1.54761e+07 muA
** NormalTransistorNmos: 1.54761e+07 muA
** NormalTransistorNmos: 4.96983e+08 muA
** NormalTransistorNmos: 4.96982e+08 muA
** NormalTransistorPmos: -4.96982e+08 muA
** NormalTransistorPmos: -4.96983e+08 muA
** DiodeTransistorNmos: 4.70111e+07 muA
** NormalTransistorNmos: 4.70111e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.16409e+07 muA
** DiodeTransistorPmos: -6.09199e+07 muA


** Expected Voltages: 
** ibias: 1.18001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.16501  V
** outInputVoltageBiasXXnXX1: 1.13601  V
** outSourceVoltageBiasXXnXX1: 0.568001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX0: 3.93701  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.87201  V
** innerTransistorStack1Load1: 4.43601  V
** innerTransistorStack2Load1: 4.43601  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.470001  V
** innerTransconductance: 4.72901  V
** inner: 0.568001  V


.END