** Name: two_stage_single_output_op_amp_44_9

.MACRO two_stage_single_output_op_amp_44_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=28e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=254e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=142e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=112e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=28e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=254e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=142e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=36e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=36e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=7e-6 W=600e-6
mMainBias17 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=595e-6
mMainBias18 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=139e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=98e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=222e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_44_9

** Expected Performance Values: 
** Gain: 118 dB
** Power consumption: 3.59001 mW
** Area: 14870 (mu_m)^2
** Transit frequency: 3.05701 MHz
** Transit frequency with error factor: 3.05699 MHz
** Slew rate: 9.77562 V/mu_s
** Phase margin: 60.7336°
** CMRR: 136 dB
** VoutMax: 4.25 V
** VoutMin: 0.710001 V
** VcmMax: 3.64001 V
** VcmMin: -0.319999 V


** Expected Currents: 
** NormalTransistorPmos: -5.33309e+07 muA
** NormalTransistorPmos: -1.23819e+07 muA
** NormalTransistorNmos: 4.47591e+07 muA
** NormalTransistorNmos: 7.18101e+07 muA
** NormalTransistorNmos: 4.47591e+07 muA
** NormalTransistorNmos: 7.18101e+07 muA
** NormalTransistorPmos: -4.47599e+07 muA
** NormalTransistorPmos: -4.47599e+07 muA
** DiodeTransistorPmos: -4.47599e+07 muA
** NormalTransistorPmos: -5.41029e+07 muA
** NormalTransistorPmos: -2.70519e+07 muA
** NormalTransistorPmos: -2.70519e+07 muA
** NormalTransistorNmos: 4.88663e+08 muA
** DiodeTransistorNmos: 4.88662e+08 muA
** NormalTransistorPmos: -4.88662e+08 muA
** DiodeTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 5.33301e+07 muA
** DiodeTransistorNmos: 1.23811e+07 muA
** DiodeTransistorNmos: 1.23801e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11101  V
** inputVoltageBiasXXnXX2: 1.20101  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.646001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.03601  V
** out1: 3.32201  V
** sourceGCC1: 0.646001  V
** sourceGCC2: 0.646001  V
** sourceTransconductance: 3.67701  V
** inner: 0.556001  V


.END