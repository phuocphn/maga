** Name: two_stage_single_output_op_amp_79_3

.MACRO two_stage_single_output_op_amp_79_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=147e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=562e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=12e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=93e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=45e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=29e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=51e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=365e-6
mFoldedCascodeFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=45e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=42e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=365e-6
mSecondStage1StageBias18 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=383e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=42e-6
mMainBias20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=544e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=109e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_79_3

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 5.49901 mW
** Area: 13177 (mu_m)^2
** Transit frequency: 4.31701 MHz
** Transit frequency with error factor: 4.31671 MHz
** Slew rate: 3.79074 V/mu_s
** Phase margin: 65.8902°
** CMRR: 149 dB
** VoutMax: 3.97001 V
** VoutMin: 0.310001 V
** VcmMax: 5.17001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorPmos: -5.51549e+08 muA
** NormalTransistorPmos: -1.10511e+08 muA
** NormalTransistorPmos: -1.71549e+07 muA
** NormalTransistorPmos: -2.63599e+07 muA
** NormalTransistorPmos: -1.71549e+07 muA
** NormalTransistorPmos: -2.63599e+07 muA
** NormalTransistorNmos: 1.71541e+07 muA
** NormalTransistorNmos: 1.71531e+07 muA
** NormalTransistorNmos: 1.71541e+07 muA
** NormalTransistorNmos: 1.71531e+07 muA
** NormalTransistorNmos: 1.84111e+07 muA
** NormalTransistorNmos: 1.84101e+07 muA
** NormalTransistorNmos: 9.20601e+06 muA
** NormalTransistorNmos: 9.20601e+06 muA
** NormalTransistorNmos: 3.65113e+08 muA
** NormalTransistorPmos: -3.65112e+08 muA
** NormalTransistorPmos: -3.65113e+08 muA
** DiodeTransistorNmos: 5.5155e+08 muA
** DiodeTransistorNmos: 1.10512e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.41801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.714001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.919001  V
** outVoltageBiasXXnXX2: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.354001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.13301  V
** sourceGCC2: 4.13301  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 4.21201  V


.END