** Name: two_stage_single_output_op_amp_122_12

.MACRO two_stage_single_output_op_amp_122_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=9e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=562e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=349e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=583e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=40e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=22e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=7e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=7e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=7e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=562e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mSecondStage1StageBias13 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=583e-6
mTelescopicFirstStageLoad14 outFirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=7e-6
mMainBias15 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=142e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=580e-6
mTelescopicFirstStageStageBias17 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=349e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=49e-6
mTelescopicFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=49e-6
mTelescopicFirstStageLoad20 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=11e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=316e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=597e-6
mTelescopicFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=11e-6
mMainBias24 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=37e-6
mMainBias25 outVoltageBiasXXnXX3 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=21e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_122_12

** Expected Performance Values: 
** Gain: 188 dB
** Power consumption: 9.43101 mW
** Area: 14297 (mu_m)^2
** Transit frequency: 3.14001 MHz
** Transit frequency with error factor: 3.14027 MHz
** Slew rate: 25.8875 V/mu_s
** Phase margin: 71.6198°
** CMRR: 129 dB
** VoutMax: 4.17001 V
** VoutMin: 0.730001 V
** VcmMax: 4.99001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 1.59324e+08 muA
** NormalTransistorNmos: 6.41953e+08 muA
** NormalTransistorPmos: -2.676e+08 muA
** NormalTransistorPmos: -1.52844e+08 muA
** NormalTransistorNmos: 6.66701e+06 muA
** NormalTransistorNmos: 6.66701e+06 muA
** NormalTransistorPmos: -6.66799e+06 muA
** NormalTransistorPmos: -6.66899e+06 muA
** NormalTransistorPmos: -6.66799e+06 muA
** NormalTransistorPmos: -6.66899e+06 muA
** NormalTransistorNmos: 1.6618e+08 muA
** DiodeTransistorNmos: 1.6618e+08 muA
** NormalTransistorNmos: 6.66701e+06 muA
** NormalTransistorNmos: 6.66701e+06 muA
** NormalTransistorNmos: 6.41172e+08 muA
** DiodeTransistorNmos: 6.41173e+08 muA
** NormalTransistorPmos: -6.41171e+08 muA
** NormalTransistorPmos: -6.41172e+08 muA
** DiodeTransistorNmos: 2.67601e+08 muA
** NormalTransistorNmos: 2.67601e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 1.52845e+08 muA
** DiodeTransistorPmos: -1.59323e+08 muA
** DiodeTransistorPmos: -6.41952e+08 muA


** Expected Voltages: 
** ibias: 1.13301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.85301  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.567001  V
** outVoltageBiasXXnXX3: 2.65001  V
** outVoltageBiasXXpXX0: 2.74501  V
** outVoltageBiasXXpXX1: 3.60901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.35701  V
** innerTransistorStack2Load2: 4.35701  V
** out1: 4.17301  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.41701  V
** inner: 0.555001  V
** inner: 0.566001  V


.END