** Name: two_stage_single_output_op_amp_8_12

.MACRO two_stage_single_output_op_amp_8_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=16e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=164e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=255e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=174e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=40e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=17e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=164e-6
mMainBias10 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=72e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=255e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=17e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=196e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=578e-6
mSecondStage1Transconductor15 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=594e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=174e-6
mMainBias17 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=406e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10e-12
.EOM two_stage_single_output_op_amp_8_12

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 8.41801 mW
** Area: 10056 (mu_m)^2
** Transit frequency: 8.22601 MHz
** Transit frequency with error factor: 8.1807 MHz
** Slew rate: 22.9288 V/mu_s
** Phase margin: 60.1606°
** CMRR: 85 dB
** negPSRR: 113 dB
** posPSRR: 83 dB
** VoutMax: 4.49001 V
** VoutMin: 0.760001 V
** VcmMax: 4.60001 V
** VcmMin: 1.30001 V


** Expected Currents: 
** NormalTransistorNmos: 4.41671e+07 muA
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorPmos: -4.40409e+08 muA
** DiodeTransistorPmos: -1.87519e+08 muA
** NormalTransistorPmos: -1.87519e+08 muA
** NormalTransistorNmos: 3.75038e+08 muA
** NormalTransistorNmos: 1.8752e+08 muA
** NormalTransistorNmos: 1.8752e+08 muA
** NormalTransistorNmos: 6.92124e+08 muA
** DiodeTransistorNmos: 6.92123e+08 muA
** NormalTransistorPmos: -6.92123e+08 muA
** NormalTransistorPmos: -6.92122e+08 muA
** DiodeTransistorNmos: 4.4041e+08 muA
** NormalTransistorNmos: 4.4041e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.41679e+07 muA
** DiodeTransistorPmos: -1.21839e+08 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.69401  V
** out: 2.5  V
** outFirstStage: 4.17701  V
** outInputVoltageBiasXXnXX1: 1.16801  V
** outSourceVoltageBiasXXnXX1: 0.584001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.19001  V
** sourceTransconductance: 1.37001  V
** innerTransconductance: 4.50501  V
** inner: 0.584001  V


.END