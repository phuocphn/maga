** Name: two_stage_single_output_op_amp_205_7

.MACRO two_stage_single_output_op_amp_205_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=28e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=28e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=56e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=10e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=28e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=22e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=45e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=383e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=28e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=22e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=136e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=136e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=434e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=200e-6
mSimpleFirstStageLoad18 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=434e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=37e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_205_7

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 6.96401 mW
** Area: 9069 (mu_m)^2
** Transit frequency: 4.78101 MHz
** Transit frequency with error factor: 4.77818 MHz
** Slew rate: 4.50601 V/mu_s
** Phase margin: 61.8795°
** CMRR: 119 dB
** VoutMax: 4.25 V
** VoutMin: 0.25 V
** VcmMax: 4.58001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorPmos: -3.70969e+07 muA
** NormalTransistorPmos: -4.97649e+07 muA
** DiodeTransistorNmos: 1.24855e+08 muA
** NormalTransistorNmos: 1.24856e+08 muA
** NormalTransistorNmos: 1.24857e+08 muA
** DiodeTransistorNmos: 1.24856e+08 muA
** NormalTransistorPmos: -1.3533e+08 muA
** NormalTransistorPmos: -1.35331e+08 muA
** NormalTransistorPmos: -1.35332e+08 muA
** NormalTransistorPmos: -1.35331e+08 muA
** NormalTransistorNmos: 2.09521e+07 muA
** NormalTransistorNmos: 2.09531e+07 muA
** NormalTransistorNmos: 1.04761e+07 muA
** NormalTransistorNmos: 1.04761e+07 muA
** NormalTransistorNmos: 1.01534e+09 muA
** NormalTransistorPmos: -1.01533e+09 muA
** DiodeTransistorNmos: 3.70961e+07 muA
** DiodeTransistorNmos: 4.97641e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.12201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 3.90901  V
** outVoltageBiasXXnXX1: 1.01501  V
** outVoltageBiasXXnXX2: 0.655001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.13401  V
** innerStageBias: 0.428001  V
** innerTransistorStack1Load1: 1.13501  V
** innerTransistorStack1Load2: 3.98001  V
** innerTransistorStack2Load2: 3.98001  V
** out1: 2.10401  V
** sourceTransconductance: 1.94501  V


.END