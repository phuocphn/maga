** Name: two_stage_single_output_op_amp_73_7

.MACRO two_stage_single_output_op_amp_73_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=139e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=22e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=49e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=139e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=11e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=11e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=94e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=587e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=5e-6 W=137e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=171e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=115e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=115e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=336e-6
mFoldedCascodeFirstStageLoad17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=171e-6
mMainBias18 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=59e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=42e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.70001e-12
.EOM two_stage_single_output_op_amp_73_7

** Expected Performance Values: 
** Gain: 115 dB
** Power consumption: 7.46001 mW
** Area: 7982 (mu_m)^2
** Transit frequency: 5.68001 MHz
** Transit frequency with error factor: 5.67982 MHz
** Slew rate: 10.2444 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 4.25 V
** VoutMin: 0.340001 V
** VcmMax: 5.17001 V
** VcmMin: 1.73001 V


** Expected Currents: 
** NormalTransistorPmos: -5.98179e+07 muA
** NormalTransistorPmos: -4.18829e+07 muA
** NormalTransistorPmos: -6.94489e+07 muA
** NormalTransistorPmos: -1.16595e+08 muA
** NormalTransistorPmos: -6.94489e+07 muA
** NormalTransistorPmos: -1.16595e+08 muA
** NormalTransistorNmos: 6.94481e+07 muA
** NormalTransistorNmos: 6.94481e+07 muA
** DiodeTransistorNmos: 6.94481e+07 muA
** NormalTransistorNmos: 9.42911e+07 muA
** NormalTransistorNmos: 9.42901e+07 muA
** NormalTransistorNmos: 4.71461e+07 muA
** NormalTransistorNmos: 4.71461e+07 muA
** NormalTransistorNmos: 1.13719e+09 muA
** NormalTransistorPmos: -1.13718e+09 muA
** DiodeTransistorNmos: 5.98171e+07 muA
** DiodeTransistorNmos: 4.18821e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.13001  V
** outVoltageBiasXXnXX2: 0.742001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.608001  V
** innerStageBias: 0.537001  V
** out1: 1.18601  V
** sourceGCC1: 4.11201  V
** sourceGCC2: 4.11201  V
** sourceTransconductance: 1.70401  V


.END