** Name: two_stage_single_output_op_amp_116_12

.MACRO two_stage_single_output_op_amp_116_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=5e-6 W=8e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=10e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=117e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=451e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=51e-6
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=10e-6 W=129e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=43e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=15e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=60e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=60e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias13 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=42e-6
mSecondStage1StageBias15 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=5e-6 W=451e-6
mTelescopicFirstStageLoad16 outFirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=15e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=271e-6
mTelescopicFirstStageStageBias18 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=117e-6
mTelescopicFirstStageLoad19 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=10e-6 W=129e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=528e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=598e-6
mTelescopicFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=3e-6 W=20e-6
mMainBias23 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=16e-6
mMainBias24 outVoltageBiasXXnXX3 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=163e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.80001e-12
.EOM two_stage_single_output_op_amp_116_12

** Expected Performance Values: 
** Gain: 181 dB
** Power consumption: 5.98701 mW
** Area: 14991 (mu_m)^2
** Transit frequency: 3.09001 MHz
** Transit frequency with error factor: 3.09003 MHz
** Slew rate: 18.4451 V/mu_s
** Phase margin: 60.1606°
** CMRR: 127 dB
** VoutMax: 4.08001 V
** VoutMin: 0.940001 V
** VcmMax: 4.09001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 5.17041e+07 muA
** NormalTransistorNmos: 3.38446e+08 muA
** NormalTransistorPmos: -1.92399e+07 muA
** NormalTransistorPmos: -1.94271e+08 muA
** NormalTransistorNmos: 1.42851e+07 muA
** NormalTransistorNmos: 1.42851e+07 muA
** NormalTransistorPmos: -1.42859e+07 muA
** NormalTransistorPmos: -1.42859e+07 muA
** DiodeTransistorPmos: -1.42859e+07 muA
** NormalTransistorNmos: 2.22843e+08 muA
** DiodeTransistorNmos: 2.22843e+08 muA
** NormalTransistorNmos: 1.42851e+07 muA
** NormalTransistorNmos: 1.42851e+07 muA
** NormalTransistorNmos: 5.55202e+08 muA
** DiodeTransistorNmos: 5.55203e+08 muA
** NormalTransistorPmos: -5.55201e+08 muA
** NormalTransistorPmos: -5.55202e+08 muA
** DiodeTransistorNmos: 1.92391e+07 muA
** NormalTransistorNmos: 1.92381e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 1.94272e+08 muA
** DiodeTransistorPmos: -5.17049e+07 muA
** DiodeTransistorPmos: -3.38445e+08 muA


** Expected Voltages: 
** ibias: 1.35001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.06901  V
** out: 2.5  V
** outFirstStage: 3.83901  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.676001  V
** outVoltageBiasXXnXX3: 2.65001  V
** outVoltageBiasXXpXX1: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.18601  V
** out1: 3.27501  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 2.82101  V
** inner: 0.554001  V
** inner: 0.672001  V


.END