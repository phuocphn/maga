** Name: two_stage_single_output_op_amp_130_3

.MACRO two_stage_single_output_op_amp_130_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=12e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=15e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=320e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=320e-6
mSimpleFirstStageLoad8 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=298e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=136e-6
mSimpleFirstStageLoad10 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=298e-6
mMainBias11 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=115e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=106e-6
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=89e-6
mSimpleFirstStageLoad14 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=155e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=596e-6
mSecondStage1StageBias17 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=494e-6
mSimpleFirstStageLoad18 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=19e-6
mSimpleFirstStageTransconductor19 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=89e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.10001e-12
.EOM two_stage_single_output_op_amp_130_3

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 7.25301 mW
** Area: 8078 (mu_m)^2
** Transit frequency: 9.08301 MHz
** Transit frequency with error factor: 9.05068 MHz
** Slew rate: 34.7119 V/mu_s
** Phase margin: 60.1606°
** CMRR: 77 dB
** VoutMax: 4.27001 V
** VoutMin: 0.390001 V
** VcmMax: 3.40001 V
** VcmMin: -0.25 V


** Expected Currents: 
** NormalTransistorNmos: 7.61491e+07 muA
** NormalTransistorNmos: 6.98781e+07 muA
** NormalTransistorPmos: -9.64569e+07 muA
** NormalTransistorPmos: -9.64559e+07 muA
** DiodeTransistorPmos: -9.64569e+07 muA
** NormalTransistorNmos: 2.09413e+08 muA
** NormalTransistorNmos: 2.09412e+08 muA
** NormalTransistorNmos: 2.09412e+08 muA
** NormalTransistorNmos: 2.09412e+08 muA
** NormalTransistorPmos: -2.25912e+08 muA
** NormalTransistorPmos: -1.12955e+08 muA
** NormalTransistorPmos: -1.12955e+08 muA
** NormalTransistorNmos: 8.75765e+08 muA
** NormalTransistorPmos: -8.75764e+08 muA
** NormalTransistorPmos: -8.75765e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.61499e+07 muA
** DiodeTransistorPmos: -6.98789e+07 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.797001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.14901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.571001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.571001  V
** out1: 2.37201  V
** sourceTransconductance: 3.81401  V
** innerStageBias: 4.69401  V


.END