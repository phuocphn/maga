** Name: two_stage_single_output_op_amp_15_4

.MACRO two_stage_single_output_op_amp_15_4 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=157e-6
mSecondStage1StageBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=59e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=13e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor5 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=318e-6
mSecondStage1Transconductor6 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=455e-6
mSimpleFirstStageLoad7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=157e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=120e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=498e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=79e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=495e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=498e-6
mMainBias14 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=266e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.60001e-12
.EOM two_stage_single_output_op_amp_15_4

** Expected Performance Values: 
** Gain: 144 dB
** Power consumption: 5.09801 mW
** Area: 10475 (mu_m)^2
** Transit frequency: 14.1631 MHz
** Transit frequency with error factor: 14.1403 MHz
** Slew rate: 18.0215 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 99 dB
** posPSRR: 114 dB
** VoutMax: 3.94001 V
** VoutMin: 0.330001 V
** VcmMax: 3.14001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorPmos: -2.6969e+08 muA
** DiodeTransistorNmos: 6.08321e+07 muA
** NormalTransistorNmos: 6.08321e+07 muA
** NormalTransistorPmos: -1.21665e+08 muA
** NormalTransistorPmos: -1.21664e+08 muA
** NormalTransistorPmos: -6.08329e+07 muA
** NormalTransistorPmos: -6.08329e+07 muA
** NormalTransistorNmos: 6.08328e+08 muA
** NormalTransistorNmos: 6.08327e+08 muA
** NormalTransistorPmos: -6.08327e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** DiodeTransistorNmos: 2.69691e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.42701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.732001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.28401  V
** out1: 0.556001  V
** sourceTransconductance: 3.26601  V
** innerStageBias: 4.25201  V
** innerTransconductance: 0.150001  V


.END