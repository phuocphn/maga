** Name: two_stage_single_output_op_amp_52_8

.MACRO two_stage_single_output_op_amp_52_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=75e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=13e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=75e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=42e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=42e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=314e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=332e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=40e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=166e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=91e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=91e-6
mMainBias16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=130e-6
mMainBias17 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=86e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=530e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=166e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.20001e-12
.EOM two_stage_single_output_op_amp_52_8

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 6.65901 mW
** Area: 6980 (mu_m)^2
** Transit frequency: 4.47801 MHz
** Transit frequency with error factor: 4.47781 MHz
** Slew rate: 4.64332 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.540001 V
** VcmMax: 5.15001 V
** VcmMin: 0.810001 V


** Expected Currents: 
** NormalTransistorPmos: -7.62869e+07 muA
** NormalTransistorPmos: -5.07929e+07 muA
** NormalTransistorPmos: -3.37089e+07 muA
** NormalTransistorPmos: -5.42449e+07 muA
** NormalTransistorPmos: -3.37089e+07 muA
** NormalTransistorPmos: -5.42449e+07 muA
** DiodeTransistorNmos: 3.37081e+07 muA
** NormalTransistorNmos: 3.37081e+07 muA
** NormalTransistorNmos: 3.37081e+07 muA
** NormalTransistorNmos: 4.10691e+07 muA
** NormalTransistorNmos: 2.05351e+07 muA
** NormalTransistorNmos: 2.05351e+07 muA
** NormalTransistorNmos: 1.07627e+09 muA
** NormalTransistorNmos: 1.07626e+09 muA
** NormalTransistorPmos: -1.07626e+09 muA
** DiodeTransistorNmos: 7.62861e+07 muA
** DiodeTransistorNmos: 5.07921e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.14401  V
** inputVoltageBiasXXnXX2: 0.606001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.17901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.566001  V
** out1: 0.568001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.89301  V
** innerStageBias: 0.401001  V


.END