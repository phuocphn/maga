** Name: one_stage_single_output_op_amp64

.MACRO one_stage_single_output_op_amp64 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=300e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=160e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=10e-6 W=122e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=10e-6 W=86e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=12e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=124e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=50e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=50e-6
mFoldedCascodeFirstStageLoad10 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=10e-6 W=122e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=373e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=373e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=124e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mMainBias16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=477e-6
mFoldedCascodeFirstStageLoad17 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=10e-6 W=86e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp64

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 3.33701 mW
** Area: 11442 (mu_m)^2
** Transit frequency: 3.83401 MHz
** Transit frequency with error factor: 3.83372 MHz
** Slew rate: 3.66188 V/mu_s
** Phase margin: 88.8085°
** CMRR: 125 dB
** VoutMax: 3.17001 V
** VoutMin: 0.840001 V
** VcmMax: 3.04001 V
** VcmMin: -0.319999 V


** Expected Currents: 
** NormalTransistorPmos: -3.9592e+08 muA
** NormalTransistorNmos: 7.33541e+07 muA
** NormalTransistorNmos: 1.25752e+08 muA
** NormalTransistorNmos: 7.33501e+07 muA
** NormalTransistorNmos: 1.25746e+08 muA
** DiodeTransistorPmos: -7.33529e+07 muA
** DiodeTransistorPmos: -7.33519e+07 muA
** NormalTransistorPmos: -7.33509e+07 muA
** NormalTransistorPmos: -7.33519e+07 muA
** NormalTransistorPmos: -1.0479e+08 muA
** DiodeTransistorPmos: -1.04789e+08 muA
** NormalTransistorPmos: -5.23959e+07 muA
** NormalTransistorPmos: -5.23959e+07 muA
** DiodeTransistorNmos: 3.95921e+08 muA
** DiodeTransistorNmos: 3.95922e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.25701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.22901  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.648001  V
** outSourceVoltageBiasXXpXX1: 4.13001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 3.85401  V
** innerTransistorStack2Load2: 3.84801  V
** out1: 2.59601  V
** sourceGCC1: 0.632001  V
** sourceGCC2: 0.632001  V
** sourceTransconductance: 3.28101  V
** inner: 4.125  V


.END