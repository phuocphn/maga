** Name: two_stage_single_output_op_amp_2_6

.MACRO two_stage_single_output_op_amp_2_6 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=41e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSecondStage1StageBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=113e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=6e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=241e-6
mSimpleFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=41e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=294e-6
mMainBias9 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=25e-6
mSecondStage1Transconductor10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=302e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=7e-6 W=41e-6
mSimpleFirstStageTransconductor12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=176e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=7e-6 W=248e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=6e-6
mMainBias15 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=25e-6
mMainBias16 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=586e-6
mSecondStage1StageBias17 out inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=241e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=176e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_2_6

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 3.35601 mW
** Area: 14985 (mu_m)^2
** Transit frequency: 4.63501 MHz
** Transit frequency with error factor: 4.63293 MHz
** Slew rate: 4.91141 V/mu_s
** Phase margin: 71.6198°
** CMRR: 105 dB
** negPSRR: 101 dB
** posPSRR: 106 dB
** VoutMax: 3 V
** VoutMin: 0.590001 V
** VcmMax: 4.08001 V
** VcmMin: 0.140001 V


** Expected Currents: 
** NormalTransistorNmos: 1.39181e+07 muA
** NormalTransistorPmos: -2.25399e+06 muA
** NormalTransistorPmos: -5.19269e+07 muA
** NormalTransistorNmos: 1.11801e+07 muA
** NormalTransistorNmos: 1.11801e+07 muA
** DiodeTransistorNmos: 1.11801e+07 muA
** NormalTransistorPmos: -2.23619e+07 muA
** NormalTransistorPmos: -1.11809e+07 muA
** NormalTransistorPmos: -1.11809e+07 muA
** NormalTransistorNmos: 5.60654e+08 muA
** NormalTransistorNmos: 5.60653e+08 muA
** NormalTransistorPmos: -5.60653e+08 muA
** DiodeTransistorPmos: -5.60653e+08 muA
** DiodeTransistorNmos: 2.25301e+06 muA
** DiodeTransistorNmos: 5.19261e+07 muA
** DiodeTransistorPmos: -1.39189e+07 muA
** NormalTransistorPmos: -1.39199e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.568001  V
** inputVoltageBiasXXnXX1: 1  V
** inputVoltageBiasXXpXX1: 2.43601  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outSourceVoltageBiasXXpXX1: 3.71801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** out1: 1.11001  V
** sourceTransconductance: 3.23201  V
** innerTransconductance: 0.300001  V
** inner: 3.71701  V


.END