** Name: two_stage_single_output_op_amp_45_7

.MACRO two_stage_single_output_op_amp_45_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=10e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=100e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=506e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=20e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=120e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=281e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=281e-6
mMainBias9 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=26e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=420e-6
mFoldedCascodeFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=120e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=506e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=67e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=67e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=467e-6
mMainBias16 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=102e-6
mMainBias17 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=207e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=568e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.6001e-12
.EOM two_stage_single_output_op_amp_45_7

** Expected Performance Values: 
** Gain: 112 dB
** Power consumption: 11.1481 mW
** Area: 7511 (mu_m)^2
** Transit frequency: 6.76401 MHz
** Transit frequency with error factor: 6.76396 MHz
** Slew rate: 23.1947 V/mu_s
** Phase margin: 60.1606°
** CMRR: 124 dB
** VoutMax: 4.73001 V
** VoutMin: 0.150001 V
** VcmMax: 3.48001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 5.00201e+07 muA
** NormalTransistorPmos: -9.40379e+07 muA
** NormalTransistorPmos: -1.90463e+08 muA
** NormalTransistorNmos: 3.19926e+08 muA
** NormalTransistorNmos: 5.35201e+08 muA
** NormalTransistorNmos: 3.19925e+08 muA
** NormalTransistorNmos: 5.35201e+08 muA
** DiodeTransistorPmos: -3.19925e+08 muA
** NormalTransistorPmos: -3.19924e+08 muA
** NormalTransistorPmos: -3.19925e+08 muA
** NormalTransistorPmos: -4.30548e+08 muA
** NormalTransistorPmos: -2.15274e+08 muA
** NormalTransistorPmos: -2.15274e+08 muA
** NormalTransistorNmos: 8.04663e+08 muA
** NormalTransistorPmos: -8.04662e+08 muA
** DiodeTransistorNmos: 9.40371e+07 muA
** DiodeTransistorNmos: 1.90464e+08 muA
** DiodeTransistorPmos: -5.00209e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.15001  V
** inputVoltageBiasXXnXX2: 0.555001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.16101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.60401  V
** out1: 4.24701  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.79501  V


.END