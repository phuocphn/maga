** Name: two_stage_single_output_op_amp_62_12

.MACRO two_stage_single_output_op_amp_62_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=8e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=355e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=106e-6
mMainBias6 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=236e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=27e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=30e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=30e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=13e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=355e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=27e-6
mMainBias15 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=106e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=450e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=450e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=236e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=492e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias22 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=58e-6
mSecondStage1Transconductor23 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=589e-6
mFoldedCascodeFirstStageLoad24 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=350e-6
mMainBias25 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=49e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 21e-12
.EOM two_stage_single_output_op_amp_62_12

** Expected Performance Values: 
** Gain: 156 dB
** Power consumption: 11.7551 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 5.58901 MHz
** Transit frequency with error factor: 5.5892 MHz
** Slew rate: 11.3334 V/mu_s
** Phase margin: 63.5984°
** CMRR: 123 dB
** VoutMax: 4.25 V
** VoutMin: 1.60001 V
** VcmMax: 3.07001 V
** VcmMin: 0.190001 V


** Expected Currents: 
** NormalTransistorNmos: 1.42147e+08 muA
** NormalTransistorPmos: -4.96799e+07 muA
** NormalTransistorPmos: -5.87759e+07 muA
** NormalTransistorNmos: 2.39278e+08 muA
** NormalTransistorNmos: 3.58915e+08 muA
** NormalTransistorNmos: 2.39279e+08 muA
** NormalTransistorNmos: 3.58916e+08 muA
** DiodeTransistorPmos: -2.39277e+08 muA
** NormalTransistorPmos: -2.39278e+08 muA
** NormalTransistorPmos: -2.39277e+08 muA
** NormalTransistorPmos: -2.39275e+08 muA
** DiodeTransistorPmos: -2.39274e+08 muA
** NormalTransistorPmos: -1.19637e+08 muA
** NormalTransistorPmos: -1.19637e+08 muA
** NormalTransistorNmos: 1.36261e+09 muA
** DiodeTransistorNmos: 1.36261e+09 muA
** NormalTransistorPmos: -1.3626e+09 muA
** NormalTransistorPmos: -1.3626e+09 muA
** DiodeTransistorNmos: 4.96791e+07 muA
** NormalTransistorNmos: 4.96781e+07 muA
** DiodeTransistorNmos: 5.87751e+07 muA
** DiodeTransistorNmos: 5.87741e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.42146e+08 muA


** Expected Voltages: 
** ibias: 3.39601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 2.14601  V
** out: 2.5  V
** outFirstStage: 4.04401  V
** outInputVoltageBiasXXnXX1: 2.01001  V
** outSourceVoltageBiasXXnXX1: 1.00501  V
** outSourceVoltageBiasXXnXX2: 1.15401  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.44501  V
** out1: 4.08101  V
** sourceGCC1: 1.09101  V
** sourceGCC2: 1.09101  V
** sourceTransconductance: 3.38601  V
** innerTransconductance: 4.60801  V
** inner: 1.00201  V
** inner: 4.19601  V


.END