** Name: two_stage_single_output_op_amp_99_3

.MACRO two_stage_single_output_op_amp_99_3 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=75e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=29e-6
mMainBias4 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=7e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=195e-6
mTelescopicFirstStageLoad7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=75e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=26e-6
mTelescopicFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=60e-6
mTelescopicFirstStageLoad10 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=7e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=9e-6 W=279e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=9e-6 W=279e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=120e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=597e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=7e-6
mMainBias16 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=24e-6
mTelescopicFirstStageStageBias17 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=600e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16e-12
.EOM two_stage_single_output_op_amp_99_3

** Expected Performance Values: 
** Gain: 104 dB
** Power consumption: 2.17501 mW
** Area: 9279 (mu_m)^2
** Transit frequency: 2.73101 MHz
** Transit frequency with error factor: 2.72914 MHz
** Slew rate: 6.75404 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** VoutMax: 3.75 V
** VoutMin: 0.170001 V
** VcmMax: 3 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorNmos: 5.35641e+07 muA
** NormalTransistorPmos: -4.88709e+07 muA
** NormalTransistorPmos: -3.41389e+07 muA
** NormalTransistorPmos: -3.41389e+07 muA
** DiodeTransistorNmos: 3.41381e+07 muA
** NormalTransistorNmos: 3.41381e+07 muA
** NormalTransistorPmos: -1.21839e+08 muA
** NormalTransistorPmos: -1.2184e+08 muA
** NormalTransistorPmos: -3.41379e+07 muA
** NormalTransistorPmos: -3.41379e+07 muA
** NormalTransistorNmos: 2.44359e+08 muA
** NormalTransistorPmos: -2.44358e+08 muA
** NormalTransistorPmos: -2.44357e+08 muA
** DiodeTransistorNmos: 4.88701e+07 muA
** DiodeTransistorPmos: -5.35649e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.20001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.577001  V
** outSourceVoltageBiasXXpXX2: 3.96101  V
** outVoltageBiasXXnXX0: 0.625  V
** outVoltageBiasXXpXX1: 1.00801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.31101  V
** innerStageBias: 3.91401  V
** out1: 0.569001  V
** sourceGCC1: 2.95501  V
** sourceGCC2: 2.95501  V
** innerStageBias: 3.97701  V


.END