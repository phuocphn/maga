** Name: one_stage_single_output_op_amp82

.MACRO one_stage_single_output_op_amp82 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=37e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=37e-6
mMainBias3 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=92e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=19e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=37e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=56e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=56e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=92e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias12 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=50e-6
mFoldedCascodeFirstStageLoad13 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=37e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=319e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=98e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=98e-6
mFoldedCascodeFirstStageLoad17 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=319e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp82

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 2.51501 mW
** Area: 2652 (mu_m)^2
** Transit frequency: 2.99901 MHz
** Transit frequency with error factor: 2.99948 MHz
** Slew rate: 6.45014 V/mu_s
** Phase margin: 88.8085°
** CMRR: 137 dB
** VoutMax: 3.94001 V
** VoutMin: 0.810001 V
** VcmMax: 5.06001 V
** VcmMin: 1.61001 V


** Expected Currents: 
** NormalTransistorNmos: 8.28211e+07 muA
** NormalTransistorPmos: -1.29556e+08 muA
** NormalTransistorPmos: -2.05129e+08 muA
** NormalTransistorPmos: -1.29556e+08 muA
** NormalTransistorPmos: -2.05129e+08 muA
** DiodeTransistorNmos: 1.29557e+08 muA
** NormalTransistorNmos: 1.29556e+08 muA
** NormalTransistorNmos: 1.29557e+08 muA
** DiodeTransistorNmos: 1.29556e+08 muA
** NormalTransistorNmos: 1.51145e+08 muA
** DiodeTransistorNmos: 1.51146e+08 muA
** NormalTransistorNmos: 7.55721e+07 muA
** NormalTransistorNmos: 7.55721e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -8.28219e+07 muA
** DiodeTransistorPmos: -8.28209e+07 muA


** Expected Voltages: 
** ibias: 1.20501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.603001  V
** outSourceVoltageBiasXXpXX1: 4.09301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.607001  V
** innerTransistorStack2Load2: 0.608001  V
** out1: 1.21601  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.69401  V
** inner: 0.601001  V


.END