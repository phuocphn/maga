** Name: two_stage_single_output_op_amp_76_3

.MACRO two_stage_single_output_op_amp_76_3 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=27e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=41e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=62e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=12e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=27e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=87e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=87e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=62e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=41e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=482e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=79e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=84e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=54e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=54e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=584e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
mSecondStage1StageBias19 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=84e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.40001e-12
.EOM two_stage_single_output_op_amp_76_3

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 3.95301 mW
** Area: 8708 (mu_m)^2
** Transit frequency: 8.06501 MHz
** Transit frequency with error factor: 8.06483 MHz
** Slew rate: 6.24525 V/mu_s
** Phase margin: 60.1606°
** CMRR: 142 dB
** VoutMax: 3.97001 V
** VoutMin: 0.290001 V
** VcmMax: 5.17001 V
** VcmMin: 1.49001 V


** Expected Currents: 
** NormalTransistorPmos: -2.73739e+07 muA
** NormalTransistorPmos: -4.15689e+07 muA
** NormalTransistorPmos: -3.40369e+07 muA
** NormalTransistorPmos: -5.47489e+07 muA
** NormalTransistorPmos: -3.40369e+07 muA
** NormalTransistorPmos: -5.47489e+07 muA
** DiodeTransistorNmos: 3.40361e+07 muA
** NormalTransistorNmos: 3.40361e+07 muA
** NormalTransistorNmos: 3.40361e+07 muA
** NormalTransistorNmos: 4.14251e+07 muA
** DiodeTransistorNmos: 4.14241e+07 muA
** NormalTransistorNmos: 2.07131e+07 muA
** NormalTransistorNmos: 2.07131e+07 muA
** NormalTransistorNmos: 5.92106e+08 muA
** NormalTransistorPmos: -5.92105e+08 muA
** NormalTransistorPmos: -5.92104e+08 muA
** DiodeTransistorNmos: 2.73731e+07 muA
** NormalTransistorNmos: 2.73721e+07 muA
** DiodeTransistorNmos: 4.15681e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.41801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.10401  V
** out: 2.5  V
** outFirstStage: 0.699001  V
** outInputVoltageBiasXXnXX1: 1.34201  V
** outSourceVoltageBiasXXnXX1: 0.671001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.498001  V
** out1: 0.703001  V
** sourceGCC1: 4.13201  V
** sourceGCC2: 4.13201  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 4.21601  V
** inner: 0.670001  V


.END