** Name: two_stage_single_output_op_amp_30_12

.MACRO two_stage_single_output_op_amp_30_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=10e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=95e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=419e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=462e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=485e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=73e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=31e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=419e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=95e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=84e-6
mSecondStage1StageBias13 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=462e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=31e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=257e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=599e-6
mSecondStage1Transconductor17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
mSimpleFirstStageLoad18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=485e-6
mMainBias19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=64e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.5e-12
.EOM two_stage_single_output_op_amp_30_12

** Expected Performance Values: 
** Gain: 131 dB
** Power consumption: 6.03201 mW
** Area: 9512 (mu_m)^2
** Transit frequency: 6.57601 MHz
** Transit frequency with error factor: 6.53809 MHz
** Slew rate: 14.7445 V/mu_s
** Phase margin: 60.1606°
** CMRR: 87 dB
** negPSRR: 112 dB
** posPSRR: 84 dB
** VoutMax: 4.59001 V
** VoutMin: 0.710001 V
** VcmMax: 4.65001 V
** VcmMin: 1.89001 V


** Expected Currents: 
** NormalTransistorNmos: 8.40661e+07 muA
** NormalTransistorNmos: 2.53835e+08 muA
** NormalTransistorPmos: -7.40199e+07 muA
** DiodeTransistorPmos: -1.65647e+08 muA
** NormalTransistorPmos: -1.65647e+08 muA
** NormalTransistorNmos: 3.31294e+08 muA
** DiodeTransistorNmos: 3.31293e+08 muA
** NormalTransistorNmos: 1.65648e+08 muA
** NormalTransistorNmos: 1.65648e+08 muA
** NormalTransistorNmos: 4.53211e+08 muA
** DiodeTransistorNmos: 4.53212e+08 muA
** NormalTransistorPmos: -4.5321e+08 muA
** NormalTransistorPmos: -4.53211e+08 muA
** DiodeTransistorNmos: 7.40191e+07 muA
** NormalTransistorNmos: 7.40191e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -8.40669e+07 muA
** DiodeTransistorPmos: -2.53834e+08 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.18101  V
** out: 2.5  V
** outFirstStage: 4.23001  V
** outInputVoltageBiasXXnXX1: 1.14401  V
** outSourceVoltageBiasXXnXX1: 0.572001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.24001  V
** sourceTransconductance: 1.34501  V
** innerTransconductance: 4.45501  V
** inner: 0.572001  V
** inner: 0.556001  V


.END