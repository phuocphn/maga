** Name: two_stage_single_output_op_amp_117_7

.MACRO two_stage_single_output_op_amp_117_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=15e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=54e-6
mTelescopicFirstStageLoad4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=204e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=29e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=25e-6
mTelescopicFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=298e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=72e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=36e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=36e-6
mMainBias11 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=172e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=72e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=50e-6
mTelescopicFirstStageStageBias15 sourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=8e-6 W=479e-6
mTelescopicFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=204e-6
mMainBias17 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=19e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=574e-6
mTelescopicFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=227e-6
mMainBias20 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=89e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.6001e-12
.EOM two_stage_single_output_op_amp_117_7

** Expected Performance Values: 
** Gain: 150 dB
** Power consumption: 2.27001 mW
** Area: 14981 (mu_m)^2
** Transit frequency: 2.74101 MHz
** Transit frequency with error factor: 2.74123 MHz
** Slew rate: 6.10074 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 4.85001 V
** VoutMin: 0.150001 V
** VcmMax: 4.38001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 6.55201e+07 muA
** NormalTransistorPmos: -6.83279e+07 muA
** NormalTransistorPmos: -1.44289e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** DiodeTransistorPmos: -2.28569e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorNmos: 1.14041e+08 muA
** NormalTransistorNmos: 1.1404e+08 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.30864e+08 muA
** NormalTransistorPmos: -2.30863e+08 muA
** DiodeTransistorNmos: 6.83271e+07 muA
** DiodeTransistorNmos: 1.44281e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** DiodeTransistorPmos: -6.55209e+07 muA


** Expected Voltages: 
** ibias: 0.555001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.705001  V
** inputVoltageBiasXXpXX1: 3.72201  V
** out: 2.5  V
** outFirstStage: 4.28601  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 3.97301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.150001  V
** innerTransistorStack2Load2: 4.43601  V
** out1: 4.27701  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END