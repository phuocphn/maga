** Name: two_stage_single_output_op_amp_59_1

.MACRO two_stage_single_output_op_amp_59_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=12e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=22e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=94e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=94e-6
mMainBias9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=35e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=120e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=22e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=53e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=107e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=107e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=3e-6 W=90e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=541e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=4e-6 W=64e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_59_1

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 6.04201 mW
** Area: 4349 (mu_m)^2
** Transit frequency: 4.77301 MHz
** Transit frequency with error factor: 4.7734 MHz
** Slew rate: 5.26336 V/mu_s
** Phase margin: 69.328°
** CMRR: 137 dB
** VoutMax: 4.66001 V
** VoutMin: 0.570001 V
** VcmMax: 3.15001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 2.03771e+07 muA
** NormalTransistorNmos: 2.37921e+07 muA
** NormalTransistorNmos: 3.58071e+07 muA
** NormalTransistorNmos: 2.37921e+07 muA
** NormalTransistorNmos: 3.58071e+07 muA
** NormalTransistorPmos: -2.37929e+07 muA
** NormalTransistorPmos: -2.37929e+07 muA
** DiodeTransistorPmos: -2.37929e+07 muA
** NormalTransistorPmos: -2.40329e+07 muA
** NormalTransistorPmos: -2.40339e+07 muA
** NormalTransistorPmos: -1.20159e+07 muA
** NormalTransistorPmos: -1.20159e+07 muA
** NormalTransistorNmos: 1.09305e+09 muA
** NormalTransistorPmos: -1.09304e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.33339e+07 muA
** DiodeTransistorPmos: -2.03779e+07 muA


** Expected Voltages: 
** ibias: 1.18101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.976001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX2: 4.10001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 3.81701  V
** innerStageBias: 4.46101  V
** out1: 2.96401  V
** sourceGCC1: 0.522001  V
** sourceGCC2: 0.522001  V
** sourceTransconductance: 3.24101  V


.END