** Name: two_stage_single_output_op_amp_100_4

.MACRO two_stage_single_output_op_amp_100_4 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=100e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=492e-6
mSecondStage1StageBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=71e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos4 L=2e-6 W=8e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=95e-6
mTelescopicFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=368e-6
mMainBias7 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=11e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=434e-6
mSecondStage1Transconductor10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=432e-6
mTelescopicFirstStageLoad11 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=100e-6
mMainBias12 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=212e-6
mMainBias13 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=110e-6
mTelescopicFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=356e-6
mTelescopicFirstStageTransconductor15 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=174e-6
mTelescopicFirstStageTransconductor16 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=174e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=203e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=95e-6
mMainBias19 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=66e-6
mMainBias20 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=133e-6
mSecondStage1StageBias21 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=597e-6
mTelescopicFirstStageLoad22 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=356e-6
mTelescopicFirstStageStageBias23 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=368e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.8001e-12
.EOM two_stage_single_output_op_amp_100_4

** Expected Performance Values: 
** Gain: 146 dB
** Power consumption: 5.60101 mW
** Area: 14686 (mu_m)^2
** Transit frequency: 4.62901 MHz
** Transit frequency with error factor: 4.62472 MHz
** Slew rate: 10.5893 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** VoutMax: 3.68001 V
** VoutMin: 0.300001 V
** VcmMax: 3 V
** VcmMin: 0.170001 V


** Expected Currents: 
** NormalTransistorNmos: 5.76831e+07 muA
** NormalTransistorNmos: 3.00551e+07 muA
** NormalTransistorPmos: -1.33868e+08 muA
** NormalTransistorPmos: -2.70829e+08 muA
** NormalTransistorPmos: -9.72299e+07 muA
** NormalTransistorPmos: -9.72299e+07 muA
** DiodeTransistorNmos: 9.72291e+07 muA
** NormalTransistorNmos: 9.72291e+07 muA
** NormalTransistorPmos: -2.24518e+08 muA
** DiodeTransistorPmos: -2.24518e+08 muA
** NormalTransistorPmos: -9.72309e+07 muA
** NormalTransistorPmos: -9.72309e+07 muA
** NormalTransistorNmos: 4.13374e+08 muA
** NormalTransistorNmos: 4.13373e+08 muA
** NormalTransistorPmos: -4.13373e+08 muA
** NormalTransistorPmos: -4.13372e+08 muA
** DiodeTransistorNmos: 1.33869e+08 muA
** DiodeTransistorNmos: 2.7083e+08 muA
** DiodeTransistorPmos: -5.76839e+07 muA
** NormalTransistorPmos: -5.76849e+07 muA
** DiodeTransistorPmos: -3.00559e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.02201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.555001  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.35201  V
** outSourceVoltageBiasXXpXX1: 4.17601  V
** outSourceVoltageBiasXXpXX3: 3.96101  V
** outVoltageBiasXXpXX2: 2.29701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.41601  V
** out1: 0.556001  V
** sourceGCC1: 3.03501  V
** sourceGCC2: 3.03501  V
** innerStageBias: 3.86301  V
** innerTransconductance: 0.150001  V
** inner: 4.17601  V


.END