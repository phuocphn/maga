** Name: two_stage_single_output_op_amp_64_2

.MACRO two_stage_single_output_op_amp_64_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=256e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=281e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=23e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=15e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=437e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=138e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=493e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=493e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=225e-6
mSecondStage1Transconductor12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=557e-6
mFoldedCascodeFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=138e-6
mMainBias14 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=256e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=78e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=78e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=437e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=11e-6
mSecondStage1StageBias21 out ibias sourcePmos sourcePmos pmos4 L=5e-6 W=600e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=281e-6
mMainBias23 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=64e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.2001e-12
.EOM two_stage_single_output_op_amp_64_2

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 3.96901 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 2.77201 MHz
** Transit frequency with error factor: 2.77188 MHz
** Slew rate: 6.56024 V/mu_s
** Phase margin: 60.1606°
** CMRR: 130 dB
** VoutMax: 4.65001 V
** VoutMin: 0.320001 V
** VcmMax: 3.06001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 6.20601e+06 muA
** NormalTransistorPmos: -2.79759e+07 muA
** NormalTransistorPmos: -4.76899e+06 muA
** NormalTransistorNmos: 1.44989e+08 muA
** NormalTransistorNmos: 2.34747e+08 muA
** NormalTransistorNmos: 1.44989e+08 muA
** NormalTransistorNmos: 2.34747e+08 muA
** DiodeTransistorPmos: -1.44988e+08 muA
** DiodeTransistorPmos: -1.44989e+08 muA
** NormalTransistorPmos: -1.44988e+08 muA
** NormalTransistorPmos: -1.44989e+08 muA
** NormalTransistorPmos: -1.79514e+08 muA
** DiodeTransistorPmos: -1.79515e+08 muA
** NormalTransistorPmos: -8.97569e+07 muA
** NormalTransistorPmos: -8.97569e+07 muA
** NormalTransistorNmos: 2.65343e+08 muA
** NormalTransistorNmos: 2.65342e+08 muA
** NormalTransistorPmos: -2.65341e+08 muA
** DiodeTransistorNmos: 2.79751e+07 muA
** DiodeTransistorNmos: 4.76801e+06 muA
** DiodeTransistorPmos: -6.20699e+06 muA
** NormalTransistorPmos: -6.20799e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.08601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.572001  V
** outInputVoltageBiasXXpXX1: 3.56801  V
** outSourceVoltageBiasXXpXX1: 4.28401  V
** outVoltageBiasXXnXX1: 0.977001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.18301  V
** innerTransistorStack2Load2: 4.18201  V
** out1: 3.37801  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.56901  V
** innerTransconductance: 0.422001  V
** inner: 4.28401  V


.END