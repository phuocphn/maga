** Name: two_stage_single_output_op_amp_75_11

.MACRO two_stage_single_output_op_amp_75_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=84e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=76e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=44e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=84e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=76e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=76e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=42e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=579e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=46e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=67e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=31e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=133e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=136e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=136e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=399e-6
mMainBias20 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=138e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=401e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=133e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.8001e-12
.EOM two_stage_single_output_op_amp_75_11

** Expected Performance Values: 
** Gain: 177 dB
** Power consumption: 7.25901 mW
** Area: 7840 (mu_m)^2
** Transit frequency: 5.17101 MHz
** Transit frequency with error factor: 5.17118 MHz
** Slew rate: 3.63741 V/mu_s
** Phase margin: 64.1713°
** CMRR: 144 dB
** VoutMax: 4.25 V
** VoutMin: 0.440001 V
** VcmMax: 5.07001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 1.11687e+08 muA
** NormalTransistorNmos: 5.09301e+07 muA
** NormalTransistorPmos: -9.31829e+07 muA
** NormalTransistorPmos: -5.40159e+07 muA
** NormalTransistorPmos: -9.02049e+07 muA
** NormalTransistorPmos: -5.40159e+07 muA
** NormalTransistorPmos: -9.02049e+07 muA
** DiodeTransistorNmos: 5.40151e+07 muA
** NormalTransistorNmos: 5.40151e+07 muA
** NormalTransistorNmos: 5.40151e+07 muA
** NormalTransistorNmos: 7.23751e+07 muA
** NormalTransistorNmos: 7.23741e+07 muA
** NormalTransistorNmos: 3.61881e+07 muA
** NormalTransistorNmos: 3.61881e+07 muA
** NormalTransistorNmos: 1.00565e+09 muA
** NormalTransistorNmos: 1.00565e+09 muA
** NormalTransistorPmos: -1.00564e+09 muA
** NormalTransistorPmos: -1.00564e+09 muA
** DiodeTransistorNmos: 9.31821e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.11686e+08 muA
** DiodeTransistorPmos: -5.09309e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.05001  V
** out: 2.5  V
** outFirstStage: 4.05901  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.10101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.398001  V
** innerTransistorStack2Load2: 0.440001  V
** out1: 0.635001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.398001  V
** innerTransconductance: 4.62301  V


.END