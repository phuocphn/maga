** Name: two_stage_single_output_op_amp_198_7

.MACRO two_stage_single_output_op_amp_198_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=2e-6 W=9e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=91e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=97e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=10e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=91e-6
mSecondStage1StageBias12 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=386e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=9e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=97e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=131e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=131e-6
mSimpleFirstStageLoad17 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=192e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=125e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=192e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=326e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.40001e-12
.EOM two_stage_single_output_op_amp_198_7

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 9.61501 mW
** Area: 5742 (mu_m)^2
** Transit frequency: 7.14901 MHz
** Transit frequency with error factor: 7.14468 MHz
** Slew rate: 6.73793 V/mu_s
** Phase margin: 60.1606°
** CMRR: 114 dB
** VoutMax: 4.25 V
** VoutMin: 0.480001 V
** VcmMax: 4.97001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorPmos: -3.29971e+08 muA
** NormalTransistorPmos: -3.95409e+07 muA
** DiodeTransistorNmos: 1.13676e+08 muA
** DiodeTransistorNmos: 1.13675e+08 muA
** NormalTransistorNmos: 1.13674e+08 muA
** NormalTransistorNmos: 1.13675e+08 muA
** NormalTransistorPmos: -1.3215e+08 muA
** NormalTransistorPmos: -1.32149e+08 muA
** NormalTransistorPmos: -1.32148e+08 muA
** NormalTransistorPmos: -1.32149e+08 muA
** NormalTransistorNmos: 3.69491e+07 muA
** DiodeTransistorNmos: 3.69481e+07 muA
** NormalTransistorNmos: 1.84751e+07 muA
** NormalTransistorNmos: 1.84751e+07 muA
** NormalTransistorNmos: 1.26918e+09 muA
** NormalTransistorPmos: -1.26917e+09 muA
** DiodeTransistorNmos: 3.29972e+08 muA
** NormalTransistorNmos: 3.29971e+08 muA
** DiodeTransistorNmos: 3.95401e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.22601  V
** outSourceVoltageBiasXXnXX1: 0.613001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.886001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.14101  V
** innerTransistorStack1Load2: 4.15801  V
** innerTransistorStack2Load1: 1.14201  V
** innerTransistorStack2Load2: 4.15801  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 0.613001  V


.END