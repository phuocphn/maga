** Name: two_stage_single_output_op_amp_187_9

.MACRO two_stage_single_output_op_amp_187_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=17e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=6e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=253e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=32e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=72e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=21e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=95e-6
mSimpleFirstStageLoad9 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=13e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=253e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=5e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=95e-6
mSimpleFirstStageLoad15 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=459e-6
mMainBias16 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=441e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=598e-6
mSimpleFirstStageLoad18 outFirstStage ibias sourcePmos sourcePmos pmos4 L=3e-6 W=459e-6
mMainBias19 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=171e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.1001e-12
.EOM two_stage_single_output_op_amp_187_9

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 6.22501 mW
** Area: 13472 (mu_m)^2
** Transit frequency: 3.79801 MHz
** Transit frequency with error factor: 3.78843 MHz
** Slew rate: 3.57918 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** VoutMax: 4.25 V
** VoutMin: 1.46001 V
** VcmMax: 5.25 V
** VcmMin: 1.30001 V


** Expected Currents: 
** NormalTransistorPmos: -2.40199e+07 muA
** NormalTransistorPmos: -6.09509e+07 muA
** NormalTransistorNmos: 4.39621e+07 muA
** NormalTransistorNmos: 4.39631e+07 muA
** DiodeTransistorNmos: 4.39621e+07 muA
** NormalTransistorPmos: -6.40679e+07 muA
** NormalTransistorPmos: -6.40679e+07 muA
** NormalTransistorNmos: 4.02091e+07 muA
** NormalTransistorNmos: 4.02081e+07 muA
** NormalTransistorNmos: 2.01051e+07 muA
** NormalTransistorNmos: 2.01051e+07 muA
** NormalTransistorNmos: 1.01196e+09 muA
** DiodeTransistorNmos: 1.01196e+09 muA
** NormalTransistorPmos: -1.01195e+09 muA
** DiodeTransistorNmos: 2.40191e+07 muA
** NormalTransistorNmos: 2.40181e+07 muA
** DiodeTransistorNmos: 6.09501e+07 muA
** DiodeTransistorNmos: 6.09491e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.16501  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.87001  V
** outSourceVoltageBiasXXnXX1: 0.935001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.568001  V
** innerTransistorStack2Load1: 1.12901  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 0.930001  V


.END