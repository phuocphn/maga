** Name: two_stage_single_output_op_amp_40_8

.MACRO two_stage_single_output_op_amp_40_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=11e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=25e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=99e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=48e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=48e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=417e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=51e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=99e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=25e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=182e-6
mSecondStage1StageBias13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=222e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=51e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=48e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=470e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=48e-6
mMainBias18 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=34e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_40_8

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 2.89701 mW
** Area: 7370 (mu_m)^2
** Transit frequency: 4.46801 MHz
** Transit frequency with error factor: 4.46504 MHz
** Slew rate: 4.2106 V/mu_s
** Phase margin: 60.1606°
** CMRR: 110 dB
** negPSRR: 109 dB
** posPSRR: 102 dB
** VoutMax: 4.69001 V
** VoutMin: 0.810001 V
** VcmMax: 3.98001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorNmos: 1.20587e+08 muA
** NormalTransistorPmos: -9.69999e+06 muA
** DiodeTransistorPmos: -1.94289e+07 muA
** NormalTransistorPmos: -1.94299e+07 muA
** NormalTransistorPmos: -1.94289e+07 muA
** DiodeTransistorPmos: -1.94299e+07 muA
** NormalTransistorNmos: 3.88551e+07 muA
** DiodeTransistorNmos: 3.88541e+07 muA
** NormalTransistorNmos: 1.94281e+07 muA
** NormalTransistorNmos: 1.94281e+07 muA
** NormalTransistorNmos: 4.00319e+08 muA
** NormalTransistorNmos: 4.00318e+08 muA
** NormalTransistorPmos: -4.00318e+08 muA
** DiodeTransistorNmos: 9.69901e+06 muA
** NormalTransistorNmos: 9.69901e+06 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.20586e+08 muA


** Expected Voltages: 
** ibias: 1.14201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.25701  V
** out: 2.5  V
** outFirstStage: 4.12601  V
** outInputVoltageBiasXXnXX1: 1.17001  V
** outSourceVoltageBiasXXnXX1: 0.585001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.28601  V
** innerTransistorStack1Load1: 4.28601  V
** out1: 3.57201  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.483001  V
** inner: 0.585001  V


.END