** Name: two_stage_single_output_op_amp_82_11

.MACRO two_stage_single_output_op_amp_82_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=5e-6 W=31e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=31e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=8e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=74e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias7 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=547e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=77e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=5e-6 W=31e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=35e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=35e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=17e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=556e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=74e-6
mMainBias15 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=202e-6
mSecondStage1StageBias16 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=582e-6
mFoldedCascodeFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=31e-6
mMainBias18 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=398e-6
mFoldedCascodeFirstStageLoad19 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=84e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=91e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=91e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=371e-6
mSecondStage1Transconductor23 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=365e-6
mFoldedCascodeFirstStageLoad24 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=84e-6
mMainBias25 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=268e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_82_11

** Expected Performance Values: 
** Gain: 177 dB
** Power consumption: 6.58601 mW
** Area: 13726 (mu_m)^2
** Transit frequency: 5.20201 MHz
** Transit frequency with error factor: 5.20155 MHz
** Slew rate: 4.90231 V/mu_s
** Phase margin: 63.5984°
** CMRR: 147 dB
** VoutMax: 4.30001 V
** VoutMin: 0.710001 V
** VcmMax: 5.03001 V
** VcmMin: 1.46001 V


** Expected Currents: 
** NormalTransistorNmos: 3.90906e+08 muA
** NormalTransistorNmos: 1.98159e+08 muA
** NormalTransistorPmos: -9.72909e+07 muA
** NormalTransistorPmos: -2.22229e+07 muA
** NormalTransistorPmos: -3.33329e+07 muA
** NormalTransistorPmos: -2.22269e+07 muA
** NormalTransistorPmos: -3.33389e+07 muA
** DiodeTransistorNmos: 2.22241e+07 muA
** NormalTransistorNmos: 2.22251e+07 muA
** NormalTransistorNmos: 2.22261e+07 muA
** DiodeTransistorNmos: 2.22251e+07 muA
** NormalTransistorNmos: 2.22211e+07 muA
** DiodeTransistorNmos: 2.22201e+07 muA
** NormalTransistorNmos: 1.11111e+07 muA
** NormalTransistorNmos: 1.11111e+07 muA
** NormalTransistorNmos: 5.54247e+08 muA
** NormalTransistorNmos: 5.54246e+08 muA
** NormalTransistorPmos: -5.54246e+08 muA
** NormalTransistorPmos: -5.54247e+08 muA
** DiodeTransistorNmos: 9.72901e+07 muA
** NormalTransistorNmos: 9.72891e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.90905e+08 muA
** DiodeTransistorPmos: -1.98158e+08 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.05801  V
** out: 2.5  V
** outFirstStage: 4.14601  V
** outInputVoltageBiasXXnXX1: 1.30601  V
** outSourceVoltageBiasXXnXX1: 0.653001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.609001  V
** innerTransistorStack2Load2: 0.610001  V
** out1: 1.17401  V
** sourceGCC1: 4.42201  V
** sourceGCC2: 4.42201  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.579001  V
** innerTransconductance: 4.66101  V
** inner: 0.651001  V


.END