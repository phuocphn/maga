** Name: two_stage_single_output_op_amp_48_6

.MACRO two_stage_single_output_op_amp_48_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=443e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=443e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=11e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=11e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=577e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=203e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=348e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=348e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mSecondStage1Transconductor12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=598e-6
mFoldedCascodeFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=203e-6
mMainBias14 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=443e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=142e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=142e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=23e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=577e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=3e-6 W=443e-6
mMainBias23 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=231e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.5e-12
.EOM two_stage_single_output_op_amp_48_6

** Expected Performance Values: 
** Gain: 178 dB
** Power consumption: 14.9991 mW
** Area: 10841 (mu_m)^2
** Transit frequency: 21.0791 MHz
** Transit frequency with error factor: 21.0791 MHz
** Slew rate: 30.6457 V/mu_s
** Phase margin: 60.1606°
** CMRR: 130 dB
** VoutMax: 3.70001 V
** VoutMin: 0.330001 V
** VcmMax: 3.79001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.68861e+07 muA
** NormalTransistorPmos: -2.11392e+08 muA
** NormalTransistorPmos: -2.09519e+07 muA
** NormalTransistorNmos: 3.88159e+08 muA
** NormalTransistorNmos: 6.65416e+08 muA
** NormalTransistorNmos: 3.88155e+08 muA
** NormalTransistorNmos: 6.6541e+08 muA
** DiodeTransistorPmos: -3.88156e+08 muA
** NormalTransistorPmos: -3.88155e+08 muA
** NormalTransistorPmos: -3.88154e+08 muA
** DiodeTransistorPmos: -3.88155e+08 muA
** NormalTransistorPmos: -5.5451e+08 muA
** NormalTransistorPmos: -2.77255e+08 muA
** NormalTransistorPmos: -2.77255e+08 muA
** NormalTransistorNmos: 1.38985e+09 muA
** NormalTransistorNmos: 1.38985e+09 muA
** NormalTransistorPmos: -1.38984e+09 muA
** DiodeTransistorPmos: -1.38984e+09 muA
** DiodeTransistorNmos: 2.11393e+08 muA
** DiodeTransistorNmos: 2.09511e+07 muA
** DiodeTransistorPmos: -2.68869e+07 muA
** NormalTransistorPmos: -2.68879e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.570001  V
** outInputVoltageBiasXXpXX1: 3.13601  V
** outSourceVoltageBiasXXpXX1: 4.06801  V
** outVoltageBiasXXnXX1: 0.905001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.05101  V
** innerTransistorStack1Load2: 4.04801  V
** out1: 3.10201  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.39301  V
** innerTransconductance: 0.334001  V
** inner: 4.06801  V


.END