** Name: two_stage_single_output_op_amp_50_9

.MACRO two_stage_single_output_op_amp_50_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=50e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=11e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=160e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=26e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=24e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=32e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=32e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=28e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=11e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=160e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=50e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=123e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=53e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=53e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=77e-6
mFoldedCascodeFirstStageLoad17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=123e-6
mMainBias18 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=110e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=35e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_50_9

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 4.55401 mW
** Area: 6995 (mu_m)^2
** Transit frequency: 3.39401 MHz
** Transit frequency with error factor: 3.39094 MHz
** Slew rate: 3.58274 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** VoutMax: 4.25 V
** VoutMin: 1.90001 V
** VcmMax: 5.12001 V
** VcmMin: 0.830001 V


** Expected Currents: 
** NormalTransistorPmos: -5.28349e+07 muA
** NormalTransistorPmos: -1.69539e+07 muA
** NormalTransistorPmos: -1.66509e+07 muA
** NormalTransistorPmos: -2.57199e+07 muA
** NormalTransistorPmos: -1.66509e+07 muA
** NormalTransistorPmos: -2.57199e+07 muA
** DiodeTransistorNmos: 1.66501e+07 muA
** NormalTransistorNmos: 1.66501e+07 muA
** NormalTransistorNmos: 1.81351e+07 muA
** NormalTransistorNmos: 9.06801e+06 muA
** NormalTransistorNmos: 9.06801e+06 muA
** NormalTransistorNmos: 7.69546e+08 muA
** DiodeTransistorNmos: 7.69545e+08 muA
** NormalTransistorPmos: -7.69545e+08 muA
** DiodeTransistorNmos: 5.28341e+07 muA
** NormalTransistorNmos: 5.28331e+07 muA
** DiodeTransistorNmos: 1.69531e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 2.31001  V
** outSourceVoltageBiasXXnXX1: 1.15501  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** outVoltageBiasXXnXX2: 0.652001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.582001  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.91201  V
** inner: 1.15501  V


.END