** Name: two_stage_single_output_op_amp_12_10

.MACRO two_stage_single_output_op_amp_12_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias2 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mSimpleFirstStageTransconductor3 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=136e-6
mSimpleFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=43e-6
mSecondStage1StageBias5 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=463e-6
mSimpleFirstStageTransconductor6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=136e-6
mMainBias7 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=158e-6
mSimpleFirstStageLoad8 FirstStageYinnerSourceLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=86e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=47e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=47e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=357e-6
mSecondStage1Transconductor12 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
mSimpleFirstStageLoad13 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=86e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18e-12
.EOM two_stage_single_output_op_amp_12_10

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 8.27001 mW
** Area: 4907 (mu_m)^2
** Transit frequency: 6.15701 MHz
** Transit frequency with error factor: 6.15355 MHz
** Slew rate: 5.86804 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 110 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 0.300001 V
** VcmMax: 4.90001 V
** VcmMin: 0.850001 V


** Expected Currents: 
** NormalTransistorNmos: 3.95982e+08 muA
** NormalTransistorPmos: -5.29839e+07 muA
** NormalTransistorPmos: -5.29849e+07 muA
** NormalTransistorPmos: -5.29839e+07 muA
** NormalTransistorPmos: -5.29849e+07 muA
** NormalTransistorNmos: 1.05967e+08 muA
** NormalTransistorNmos: 5.29831e+07 muA
** NormalTransistorNmos: 5.29831e+07 muA
** NormalTransistorNmos: 1.14205e+09 muA
** NormalTransistorPmos: -1.14204e+09 muA
** NormalTransistorPmos: -1.14204e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.95981e+08 muA


** Expected Voltages: 
** ibias: 0.702001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.01101  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.93501  V
** innerTransistorStack1Load1: 4.43501  V
** innerTransistorStack2Load1: 4.43501  V
** sourceTransconductance: 1.94301  V
** innerTransconductance: 4.57501  V


.END