** Name: two_stage_single_output_op_amp_65_12

.MACRO two_stage_single_output_op_amp_65_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=25e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=145e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=24e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=66e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=139e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=139e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=145e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=66e-6
mMainBias13 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=111e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=600e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=129e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=129e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=301e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=489e-6
mFoldedCascodeFirstStageTransconductor19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=489e-6
mFoldedCascodeFirstStageStageBias20 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=600e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=442e-6
mMainBias22 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=523e-6
mMainBias23 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=70e-6
mSecondStage1Transconductor24 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad25 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=301e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.3001e-12
.EOM two_stage_single_output_op_amp_65_12

** Expected Performance Values: 
** Gain: 166 dB
** Power consumption: 13.1541 mW
** Area: 14889 (mu_m)^2
** Transit frequency: 6.80601 MHz
** Transit frequency with error factor: 6.80564 MHz
** Slew rate: 14.5672 V/mu_s
** Phase margin: 61.3065°
** CMRR: 132 dB
** VoutMax: 4.25 V
** VoutMin: 1.05001 V
** VcmMax: 3.12001 V
** VcmMin: -0.379999 V


** Expected Currents: 
** NormalTransistorNmos: 3.04104e+08 muA
** NormalTransistorPmos: -2.19955e+08 muA
** NormalTransistorPmos: -2.95419e+07 muA
** NormalTransistorNmos: 2.53522e+08 muA
** NormalTransistorNmos: 3.80281e+08 muA
** NormalTransistorNmos: 2.53524e+08 muA
** NormalTransistorNmos: 3.80283e+08 muA
** NormalTransistorPmos: -2.53521e+08 muA
** NormalTransistorPmos: -2.53522e+08 muA
** NormalTransistorPmos: -2.53523e+08 muA
** NormalTransistorPmos: -2.53522e+08 muA
** NormalTransistorPmos: -2.53519e+08 muA
** NormalTransistorPmos: -2.53518e+08 muA
** NormalTransistorPmos: -1.26759e+08 muA
** NormalTransistorPmos: -1.26759e+08 muA
** NormalTransistorNmos: 1.29656e+09 muA
** DiodeTransistorNmos: 1.29656e+09 muA
** NormalTransistorPmos: -1.29655e+09 muA
** NormalTransistorPmos: -1.29656e+09 muA
** DiodeTransistorNmos: 2.19956e+08 muA
** NormalTransistorNmos: 2.19957e+08 muA
** DiodeTransistorNmos: 2.95411e+07 muA
** DiodeTransistorNmos: 2.95401e+07 muA
** DiodeTransistorPmos: -3.04103e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.45801  V
** inputVoltageBiasXXnXX2: 1.17501  V
** out: 2.5  V
** outFirstStage: 4.03201  V
** outSourceVoltageBiasXXnXX1: 0.729001  V
** outSourceVoltageBiasXXnXX2: 0.584001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40301  V
** innerTransistorStack1Load2: 4.46701  V
** innerTransistorStack2Load2: 4.46701  V
** out1: 4.10301  V
** sourceGCC1: 0.556001  V
** sourceGCC2: 0.556001  V
** sourceTransconductance: 3.40301  V
** innerTransconductance: 4.59601  V
** inner: 0.730001  V


.END