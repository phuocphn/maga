** Name: two_stage_single_output_op_amp_169_6

.MACRO two_stage_single_output_op_amp_169_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=35e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=505e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=84e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=88e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=299e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad9 FirstStageYinnerOutputLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=359e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=359e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=359e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=589e-6
mSecondStage1Transconductor13 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=591e-6
mSimpleFirstStageLoad14 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=359e-6
mMainBias15 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=177e-6
mSimpleFirstStageTransconductor16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=248e-6
mSimpleFirstStageStageBias17 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=369e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=84e-6
mSimpleFirstStageStageBias19 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=185e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=88e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=299e-6
mSimpleFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=505e-6
mSimpleFirstStageTransconductor23 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=248e-6
mMainBias24 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=76e-6
mMainBias25 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=67e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.5e-12
.EOM two_stage_single_output_op_amp_169_6

** Expected Performance Values: 
** Gain: 140 dB
** Power consumption: 14.9691 mW
** Area: 7273 (mu_m)^2
** Transit frequency: 14.8761 MHz
** Transit frequency with error factor: 14.8623 MHz
** Slew rate: 27.1565 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** VoutMax: 3.13001 V
** VoutMin: 0.300001 V
** VcmMax: 3.01001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 3.3712e+08 muA
** NormalTransistorPmos: -7.69549e+07 muA
** NormalTransistorPmos: -6.66629e+07 muA
** DiodeTransistorPmos: -4.967e+08 muA
** DiodeTransistorPmos: -4.96701e+08 muA
** NormalTransistorPmos: -4.967e+08 muA
** NormalTransistorPmos: -4.96701e+08 muA
** NormalTransistorNmos: 6.83762e+08 muA
** NormalTransistorNmos: 6.83762e+08 muA
** NormalTransistorNmos: 6.83762e+08 muA
** NormalTransistorNmos: 6.83762e+08 muA
** NormalTransistorPmos: -3.74121e+08 muA
** NormalTransistorPmos: -3.7412e+08 muA
** NormalTransistorPmos: -1.8706e+08 muA
** NormalTransistorPmos: -1.8706e+08 muA
** NormalTransistorNmos: 1.12564e+09 muA
** NormalTransistorNmos: 1.12564e+09 muA
** NormalTransistorPmos: -1.12563e+09 muA
** DiodeTransistorPmos: -1.12563e+09 muA
** DiodeTransistorNmos: 7.69541e+07 muA
** DiodeTransistorNmos: 6.66621e+07 muA
** DiodeTransistorPmos: -3.37119e+08 muA
** NormalTransistorPmos: -3.3712e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.56801  V
** outSourceVoltageBiasXXpXX1: 3.78401  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX1: 0.705001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.05901  V
** innerSourceLoad1: 3.85801  V
** innerStageBias: 4.29701  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load1: 3.85701  V
** innerTransistorStack2Load2: 0.150001  V
** sourceTransconductance: 3.35401  V
** innerTransconductance: 0.150001  V
** inner: 3.78401  V


.END