** Name: two_stage_single_output_op_amp_16_1

.MACRO two_stage_single_output_op_amp_16_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=10e-6 W=27e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=28e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=53e-6
mSimpleFirstStageLoad7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mMainBias8 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=23e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=78e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=40e-6
mMainBias11 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mMainBias12 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=10e-6 W=20e-6
mSecondStage1StageBias13 out ibias sourcePmos sourcePmos pmos4 L=10e-6 W=268e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=78e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.40001e-12
.EOM two_stage_single_output_op_amp_16_1

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 0.809001 mW
** Area: 4833 (mu_m)^2
** Transit frequency: 3.06501 MHz
** Transit frequency with error factor: 3.05918 MHz
** Slew rate: 3.60969 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 101 dB
** posPSRR: 212 dB
** VoutMax: 4.54001 V
** VoutMin: 0.150001 V
** VcmMax: 3.35001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 1.39251e+07 muA
** NormalTransistorPmos: -7.39899e+06 muA
** DiodeTransistorNmos: 9.79601e+06 muA
** NormalTransistorNmos: 9.79601e+06 muA
** NormalTransistorPmos: -1.95929e+07 muA
** DiodeTransistorPmos: -1.95939e+07 muA
** NormalTransistorPmos: -9.79699e+06 muA
** NormalTransistorPmos: -9.79699e+06 muA
** NormalTransistorNmos: 1.00963e+08 muA
** NormalTransistorPmos: -1.00962e+08 muA
** DiodeTransistorNmos: 7.39801e+06 muA
** DiodeTransistorPmos: -1.39259e+07 muA
** NormalTransistorPmos: -1.39269e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 3.97901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.613001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.54001  V
** outSourceVoltageBiasXXpXX1: 4.27001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceTransconductance: 3.25101  V
** inner: 4.27001  V


.END