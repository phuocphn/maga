** Name: two_stage_single_output_op_amp_3_1

.MACRO two_stage_single_output_op_amp_3_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=115e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=115e-6
mSecondStage1Transconductor5 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=215e-6
mSimpleFirstStageLoad6 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=36e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=30e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=237e-6
mMainBias9 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
mSecondStage1StageBias10 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=446e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=30e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_3_1

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 1.77601 mW
** Area: 2524 (mu_m)^2
** Transit frequency: 5.39701 MHz
** Transit frequency with error factor: 5.37944 MHz
** Slew rate: 8.31196 V/mu_s
** Phase margin: 65.3172°
** CMRR: 93 dB
** negPSRR: 95 dB
** posPSRR: 197 dB
** VoutMax: 4.84001 V
** VoutMin: 0.150001 V
** VcmMax: 3.56001 V
** VcmMin: 0.220001 V


** Expected Currents: 
** NormalTransistorPmos: -2.09049e+07 muA
** DiodeTransistorNmos: 5.47581e+07 muA
** NormalTransistorNmos: 5.47571e+07 muA
** NormalTransistorNmos: 5.47581e+07 muA
** NormalTransistorPmos: -1.09515e+08 muA
** NormalTransistorPmos: -5.47579e+07 muA
** NormalTransistorPmos: -5.47579e+07 muA
** NormalTransistorNmos: 2.04749e+08 muA
** NormalTransistorPmos: -2.04748e+08 muA
** DiodeTransistorNmos: 2.09041e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.788001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.77601  V


.END