** Name: two_stage_single_output_op_amp_148_12

.MACRO two_stage_single_output_op_amp_148_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=7e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=34e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=416e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=185e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=148e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=196e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=34e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=416e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=7e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=148e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=536e-6
mMainBias16 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=596e-6
mSimpleFirstStageLoad17 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=162e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=84e-6
mSimpleFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=84e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=464e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=162e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=58e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.2001e-12
.EOM two_stage_single_output_op_amp_148_12

** Expected Performance Values: 
** Gain: 140 dB
** Power consumption: 12.1171 mW
** Area: 12338 (mu_m)^2
** Transit frequency: 7.36001 MHz
** Transit frequency with error factor: 7.35637 MHz
** Slew rate: 6.9492 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** VoutMax: 4.25 V
** VoutMin: 1.18001 V
** VcmMax: 4.85001 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 3.14755e+08 muA
** NormalTransistorNmos: 3.44988e+08 muA
** NormalTransistorPmos: -1.08852e+08 muA
** DiodeTransistorNmos: 1.0246e+08 muA
** DiodeTransistorNmos: 1.02459e+08 muA
** NormalTransistorNmos: 1.02458e+08 muA
** NormalTransistorNmos: 1.02459e+08 muA
** NormalTransistorPmos: -1.59042e+08 muA
** NormalTransistorPmos: -1.59041e+08 muA
** NormalTransistorPmos: -1.5904e+08 muA
** NormalTransistorPmos: -1.59041e+08 muA
** NormalTransistorNmos: 1.13168e+08 muA
** NormalTransistorNmos: 5.65831e+07 muA
** NormalTransistorNmos: 5.65831e+07 muA
** NormalTransistorNmos: 1.32672e+09 muA
** DiodeTransistorNmos: 1.32671e+09 muA
** NormalTransistorPmos: -1.32671e+09 muA
** NormalTransistorPmos: -1.32671e+09 muA
** DiodeTransistorNmos: 1.08853e+08 muA
** NormalTransistorNmos: 1.08852e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.14754e+08 muA
** DiodeTransistorPmos: -3.44987e+08 muA


** Expected Voltages: 
** ibias: 0.571001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.03601  V
** outInputVoltageBiasXXnXX1: 1.58401  V
** outSourceVoltageBiasXXnXX1: 0.792001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.11201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.10001  V
** innerTransistorStack1Load1: 1.10401  V
** innerTransistorStack1Load2: 4.48401  V
** innerTransistorStack2Load1: 1.10501  V
** innerTransistorStack2Load2: 4.48401  V
** sourceTransconductance: 1.94401  V
** innerTransconductance: 4.60001  V
** inner: 0.789001  V


.END