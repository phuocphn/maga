** Name: two_stage_single_output_op_amp_12_7

.MACRO two_stage_single_output_op_amp_12_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mMainBias2 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mSimpleFirstStageTransconductor3 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=10e-6
mSimpleFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=15e-6
mMainBias5 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=25e-6
mSecondStage1StageBias6 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=188e-6
mSimpleFirstStageTransconductor7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=10e-6
mSimpleFirstStageLoad8 FirstStageYinnerSourceLoad1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=73e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=16e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=16e-6
mSecondStage1Transconductor11 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=178e-6
mSimpleFirstStageLoad12 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=73e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_12_7

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 2.29901 mW
** Area: 2573 (mu_m)^2
** Transit frequency: 2.55001 MHz
** Transit frequency with error factor: 2.54619 MHz
** Slew rate: 5.97382 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** negPSRR: 91 dB
** posPSRR: 87 dB
** VoutMax: 4.32001 V
** VoutMin: 0.340001 V
** VcmMax: 4.81001 V
** VcmMin: 1.12001 V


** Expected Currents: 
** NormalTransistorNmos: 5.00051e+07 muA
** NormalTransistorPmos: -1.47049e+07 muA
** NormalTransistorPmos: -1.47059e+07 muA
** NormalTransistorPmos: -1.47049e+07 muA
** NormalTransistorPmos: -1.47059e+07 muA
** NormalTransistorNmos: 2.94091e+07 muA
** NormalTransistorNmos: 1.47041e+07 muA
** NormalTransistorNmos: 1.47041e+07 muA
** NormalTransistorNmos: 3.70329e+08 muA
** NormalTransistorPmos: -3.70328e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.00059e+07 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.75701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.83601  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.72101  V


.END