** Name: two_stage_single_output_op_amp_92_9

.MACRO two_stage_single_output_op_amp_92_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=19e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=538e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=28e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=17e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=71e-6
mTelescopicFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=49e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=10e-6 W=82e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=10e-6 W=82e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=538e-6
mTelescopicFirstStageLoad12 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=49e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
mTelescopicFirstStageStageBias14 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=8e-6 W=127e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=336e-6
mTelescopicFirstStageLoad16 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=17e-6
mMainBias17 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=112e-6
mMainBias18 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=161e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.5e-12
.EOM two_stage_single_output_op_amp_92_9

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 5.70801 mW
** Area: 6032 (mu_m)^2
** Transit frequency: 6.00801 MHz
** Transit frequency with error factor: 6.00556 MHz
** Slew rate: 12.0437 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** VoutMax: 4.59001 V
** VoutMin: 0.700001 V
** VcmMax: 4.30001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorNmos: 1.54901e+07 muA
** NormalTransistorPmos: -2.49149e+07 muA
** NormalTransistorPmos: -3.52019e+07 muA
** NormalTransistorNmos: 1.56171e+07 muA
** NormalTransistorNmos: 1.56171e+07 muA
** DiodeTransistorPmos: -1.56179e+07 muA
** NormalTransistorPmos: -1.56179e+07 muA
** NormalTransistorNmos: 6.64361e+07 muA
** NormalTransistorNmos: 1.56181e+07 muA
** NormalTransistorNmos: 1.56181e+07 muA
** NormalTransistorNmos: 1.02469e+09 muA
** DiodeTransistorNmos: 1.02469e+09 muA
** NormalTransistorPmos: -1.02468e+09 muA
** DiodeTransistorNmos: 2.49141e+07 muA
** NormalTransistorNmos: 2.49131e+07 muA
** DiodeTransistorNmos: 3.52011e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.54909e+07 muA


** Expected Voltages: 
** ibias: 0.627001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.02101  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 4.27901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.04201  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.554001  V


.END