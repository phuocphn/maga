** Name: symmetrical_op_amp184

.MACRO symmetrical_op_amp184 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=68e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias4 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSymmetricalFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=73e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=37e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=68e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=86e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=35e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=86e-6
mMainBias12 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=3e-6 W=28e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=41e-6
mSymmetricalFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=8e-6 W=41e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=49e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=8e-6 W=49e-6
mSymmetricalFirstStageLoad18 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=162e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor19 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=196e-6
mSecondStage1Transconductor20 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=196e-6
mSymmetricalFirstStageLoad21 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=162e-6
mMainBias22 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=15e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp184

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 1.13601 mW
** Area: 5295 (mu_m)^2
** Transit frequency: 4.14401 MHz
** Transit frequency with error factor: 4.14389 MHz
** Slew rate: 3.97017 V/mu_s
** Phase margin: 74.4846°
** CMRR: 144 dB
** negPSRR: 120 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 0.380001 V
** VcmMax: 4.81001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 9.84701e+06 muA
** NormalTransistorNmos: 2.53821e+07 muA
** NormalTransistorPmos: -3.68839e+07 muA
** NormalTransistorPmos: -3.27609e+07 muA
** NormalTransistorPmos: -3.27619e+07 muA
** NormalTransistorPmos: -3.27609e+07 muA
** NormalTransistorPmos: -3.27619e+07 muA
** NormalTransistorNmos: 6.55191e+07 muA
** NormalTransistorNmos: 6.55181e+07 muA
** NormalTransistorNmos: 3.27601e+07 muA
** NormalTransistorNmos: 3.27601e+07 muA
** NormalTransistorNmos: 3.98001e+07 muA
** NormalTransistorNmos: 3.97991e+07 muA
** NormalTransistorPmos: -3.98009e+07 muA
** NormalTransistorPmos: -3.98009e+07 muA
** DiodeTransistorNmos: 3.98001e+07 muA
** NormalTransistorPmos: -3.98009e+07 muA
** NormalTransistorPmos: -3.98009e+07 muA
** DiodeTransistorNmos: 3.68831e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.84799e+06 muA
** DiodeTransistorPmos: -2.53829e+07 muA


** Expected Voltages: 
** ibias: 0.584001  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.624001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 0.788001  V
** outVoltageBiasXXpXX0: 3.69101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.179001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.219001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END