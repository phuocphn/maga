** Name: two_stage_single_output_op_amp_44_10

.MACRO two_stage_single_output_op_amp_44_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=23e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=298e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=572e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=13e-6
mSecondStage1StageBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=45e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=51e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=218e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=218e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=470e-6
mFoldedCascodeFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=51e-6
mMainBias11 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=388e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=572e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=103e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=103e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=258e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=225e-6
mMainBias17 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=355e-6
mMainBias18 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=452e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=381e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.7001e-12
.EOM two_stage_single_output_op_amp_44_10

** Expected Performance Values: 
** Gain: 114 dB
** Power consumption: 10.8261 mW
** Area: 11663 (mu_m)^2
** Transit frequency: 2.92201 MHz
** Transit frequency with error factor: 2.92137 MHz
** Slew rate: 10.4196 V/mu_s
** Phase margin: 60.1606°
** CMRR: 127 dB
** VoutMax: 4.25 V
** VoutMin: 0.170001 V
** VcmMax: 3.41001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorNmos: 4.56903e+08 muA
** NormalTransistorPmos: -2.74347e+08 muA
** NormalTransistorPmos: -3.48277e+08 muA
** NormalTransistorNmos: 1.54506e+08 muA
** NormalTransistorNmos: 2.55139e+08 muA
** NormalTransistorNmos: 1.54507e+08 muA
** NormalTransistorNmos: 2.5514e+08 muA
** NormalTransistorPmos: -1.54505e+08 muA
** NormalTransistorPmos: -1.54506e+08 muA
** DiodeTransistorPmos: -1.54505e+08 muA
** NormalTransistorPmos: -2.01266e+08 muA
** NormalTransistorPmos: -1.00633e+08 muA
** NormalTransistorPmos: -1.00633e+08 muA
** NormalTransistorNmos: 5.55451e+08 muA
** NormalTransistorPmos: -5.5545e+08 muA
** NormalTransistorPmos: -5.55449e+08 muA
** DiodeTransistorNmos: 2.74348e+08 muA
** DiodeTransistorNmos: 3.48278e+08 muA
** DiodeTransistorPmos: -4.56902e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.14201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.15201  V
** inputVoltageBiasXXnXX2: 0.572001  V
** out: 2.5  V
** outFirstStage: 3.91301  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.26301  V
** out1: 3.54901  V
** sourceGCC1: 0.367001  V
** sourceGCC2: 0.367001  V
** sourceTransconductance: 3.80001  V
** innerTransconductance: 4.47701  V


.END