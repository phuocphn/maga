** Name: two_stage_single_output_op_amp_12_11

.MACRO two_stage_single_output_op_amp_12_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mMainBias3 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=72e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSimpleFirstStageTransconductor5 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=113e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=46e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=512e-6
mSecondStage1StageBias8 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=590e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=113e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=19e-6
mMainBias11 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=45e-6
mSimpleFirstStageLoad12 FirstStageYinnerSourceLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=104e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=36e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=36e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=425e-6
mSecondStage1Transconductor16 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad17 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=104e-6
mMainBias18 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=264e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.9001e-12
.EOM two_stage_single_output_op_amp_12_11

** Expected Performance Values: 
** Gain: 141 dB
** Power consumption: 8.55401 mW
** Area: 10539 (mu_m)^2
** Transit frequency: 7.81301 MHz
** Transit frequency with error factor: 7.80865 MHz
** Slew rate: 7.53656 V/mu_s
** Phase margin: 60.1606°
** CMRR: 101 dB
** negPSRR: 109 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 0.700001 V
** VcmMax: 4.99001 V
** VcmMin: 0.900001 V


** Expected Currents: 
** NormalTransistorNmos: 4.65651e+07 muA
** NormalTransistorNmos: 1.11687e+08 muA
** NormalTransistorPmos: -1.7052e+08 muA
** NormalTransistorPmos: -5.63679e+07 muA
** NormalTransistorPmos: -5.63689e+07 muA
** NormalTransistorPmos: -5.63679e+07 muA
** NormalTransistorPmos: -5.63689e+07 muA
** NormalTransistorNmos: 1.12736e+08 muA
** NormalTransistorNmos: 5.63671e+07 muA
** NormalTransistorNmos: 5.63671e+07 muA
** NormalTransistorNmos: 1.25936e+09 muA
** NormalTransistorNmos: 1.25936e+09 muA
** NormalTransistorPmos: -1.25935e+09 muA
** NormalTransistorPmos: -1.25935e+09 muA
** DiodeTransistorNmos: 1.70521e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.65659e+07 muA
** DiodeTransistorPmos: -1.11686e+08 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.02701  V
** outVoltageBiasXXnXX1: 1.10101  V
** outVoltageBiasXXpXX0: 3.89601  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.01601  V
** innerTransistorStack1Load1: 4.42401  V
** innerTransistorStack2Load1: 4.42401  V
** sourceTransconductance: 1.94101  V
** innerStageBias: 0.342001  V
** innerTransconductance: 4.59101  V


.END