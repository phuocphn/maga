** Name: two_stage_single_output_op_amp_81_1

.MACRO two_stage_single_output_op_amp_81_1 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=129e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=129e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=29e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=42e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=147e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=129e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=52e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=52e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=8e-6 W=91e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=10e-6 W=472e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=9e-6 W=129e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=55e-6
mMainBias15 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=118e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=78e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=78e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.40001e-12
.EOM two_stage_single_output_op_amp_81_1

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 5.65001 mW
** Area: 14995 (mu_m)^2
** Transit frequency: 5.57801 MHz
** Transit frequency with error factor: 5.57755 MHz
** Slew rate: 4.22223 V/mu_s
** Phase margin: 60.1606°
** CMRR: 144 dB
** VoutMax: 4.70001 V
** VoutMin: 0.5 V
** VcmMax: 5.10001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 1.32261e+07 muA
** NormalTransistorNmos: 2.82321e+07 muA
** NormalTransistorPmos: -2.73009e+07 muA
** NormalTransistorPmos: -4.47999e+07 muA
** NormalTransistorPmos: -2.73009e+07 muA
** NormalTransistorPmos: -4.47999e+07 muA
** DiodeTransistorNmos: 2.73001e+07 muA
** NormalTransistorNmos: 2.73001e+07 muA
** NormalTransistorNmos: 2.73001e+07 muA
** DiodeTransistorNmos: 2.73001e+07 muA
** NormalTransistorNmos: 3.49971e+07 muA
** NormalTransistorNmos: 3.49981e+07 muA
** NormalTransistorNmos: 1.74981e+07 muA
** NormalTransistorNmos: 1.74981e+07 muA
** NormalTransistorNmos: 9.88982e+08 muA
** NormalTransistorPmos: -9.88981e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.32269e+07 muA
** DiodeTransistorPmos: -2.82329e+07 muA


** Expected Voltages: 
** ibias: 1.14001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.905001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 3.68801  V
** outVoltageBiasXXpXX2: 4.13101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerStageBias: 0.544001  V
** innerTransistorStack1Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 4.49401  V
** sourceGCC2: 4.49401  V
** sourceTransconductance: 1.94001  V


.END