** Name: two_stage_single_output_op_amp_66_12

.MACRO two_stage_single_output_op_amp_66_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=5e-6 W=16e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=51e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=292e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=23e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=533e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=68e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=41e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=41e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=292e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=68e-6
mMainBias14 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=12e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=97e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=97e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=395e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=395e-6
mFoldedCascodeFirstStageTransconductor19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=395e-6
mFoldedCascodeFirstStageStageBias20 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=533e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=536e-6
mMainBias22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=23e-6
mMainBias23 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=154e-6
mSecondStage1Transconductor24 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad25 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=395e-6
mMainBias26 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=563e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.4001e-12
.EOM two_stage_single_output_op_amp_66_12

** Expected Performance Values: 
** Gain: 161 dB
** Power consumption: 12.8891 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 6.39201 MHz
** Transit frequency with error factor: 6.39177 MHz
** Slew rate: 12.7066 V/mu_s
** Phase margin: 61.8795°
** CMRR: 126 dB
** VoutMax: 4.25 V
** VoutMin: 1.08001 V
** VcmMax: 3.01001 V
** VcmMin: 0.150001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -2.4706e+08 muA
** NormalTransistorPmos: -6.76019e+07 muA
** NormalTransistorNmos: 2.35526e+08 muA
** NormalTransistorNmos: 3.53287e+08 muA
** NormalTransistorNmos: 2.35528e+08 muA
** NormalTransistorNmos: 3.53289e+08 muA
** NormalTransistorPmos: -2.35525e+08 muA
** NormalTransistorPmos: -2.35526e+08 muA
** NormalTransistorPmos: -2.35527e+08 muA
** NormalTransistorPmos: -2.35526e+08 muA
** NormalTransistorPmos: -2.35523e+08 muA
** DiodeTransistorPmos: -2.35522e+08 muA
** NormalTransistorPmos: -1.17761e+08 muA
** NormalTransistorPmos: -1.17761e+08 muA
** NormalTransistorNmos: 1.43498e+09 muA
** DiodeTransistorNmos: 1.43497e+09 muA
** NormalTransistorPmos: -1.43497e+09 muA
** NormalTransistorPmos: -1.43497e+09 muA
** DiodeTransistorNmos: 2.47061e+08 muA
** NormalTransistorNmos: 2.47062e+08 muA
** DiodeTransistorNmos: 6.76011e+07 muA
** DiodeTransistorNmos: 6.76001e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 3.32801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 2.01801  V
** out: 2.5  V
** outFirstStage: 4.05001  V
** outInputVoltageBiasXXnXX1: 1.49001  V
** outSourceVoltageBiasXXnXX1: 0.745001  V
** outSourceVoltageBiasXXnXX2: 1.11501  V
** outSourceVoltageBiasXXpXX1: 4.16501  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.43201  V
** innerTransistorStack2Load2: 4.43201  V
** out1: 4.06801  V
** sourceGCC1: 1.15901  V
** sourceGCC2: 1.15901  V
** sourceTransconductance: 3.37901  V
** innerTransconductance: 4.61401  V
** inner: 0.746001  V
** inner: 4.16101  V


.END