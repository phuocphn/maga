** Name: two_stage_single_output_op_amp_51_6

.MACRO two_stage_single_output_op_amp_51_6 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=240e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=10e-6
mSecondStage1StageBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=7e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=42e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=135e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=42e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=240e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=16e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=223e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=265e-6
mMainBias13 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=35e-6
mSecondStage1Transconductor14 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=595e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=6e-6 W=471e-6
mMainBias16 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=364e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=587e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=320e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=320e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=42e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=135e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=587e-6
mMainBias23 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=494e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.1001e-12
.EOM two_stage_single_output_op_amp_51_6

** Expected Performance Values: 
** Gain: 162 dB
** Power consumption: 12.3091 mW
** Area: 14489 (mu_m)^2
** Transit frequency: 4.97901 MHz
** Transit frequency with error factor: 4.97941 MHz
** Slew rate: 8.80486 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 3.06001 V
** VoutMin: 0.650001 V
** VcmMax: 5.10001 V
** VcmMin: 1.05001 V


** Expected Currents: 
** NormalTransistorNmos: 3.58853e+08 muA
** NormalTransistorNmos: 3.45711e+07 muA
** NormalTransistorPmos: -3.99833e+08 muA
** NormalTransistorPmos: -1.53237e+08 muA
** NormalTransistorPmos: -2.62694e+08 muA
** NormalTransistorPmos: -1.53236e+08 muA
** NormalTransistorPmos: -2.62693e+08 muA
** NormalTransistorNmos: 1.53238e+08 muA
** NormalTransistorNmos: 1.53237e+08 muA
** DiodeTransistorNmos: 1.53238e+08 muA
** NormalTransistorNmos: 2.18914e+08 muA
** NormalTransistorNmos: 1.09457e+08 muA
** NormalTransistorNmos: 1.09457e+08 muA
** NormalTransistorNmos: 1.13326e+09 muA
** NormalTransistorNmos: 1.13326e+09 muA
** NormalTransistorPmos: -1.13325e+09 muA
** DiodeTransistorPmos: -1.13325e+09 muA
** DiodeTransistorNmos: 3.99834e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.58852e+08 muA
** NormalTransistorPmos: -3.58851e+08 muA
** DiodeTransistorPmos: -3.45719e+07 muA
** DiodeTransistorPmos: -3.45709e+07 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.82301  V
** out: 2.5  V
** outFirstStage: 0.907001  V
** outInputVoltageBiasXXpXX1: 2.49601  V
** outSourceVoltageBiasXXpXX1: 3.74801  V
** outSourceVoltageBiasXXpXX2: 4.13401  V
** outVoltageBiasXXnXX1: 1.05701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** out1: 1.11201  V
** sourceGCC1: 3.55801  V
** sourceGCC2: 3.55801  V
** sourceTransconductance: 1.69101  V
** innerTransconductance: 0.502001  V
** inner: 3.74901  V


.END