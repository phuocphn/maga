** Name: two_stage_single_output_op_amp_37_9

.MACRO two_stage_single_output_op_amp_37_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=7e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=411e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=5e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=7e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=19e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=19e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=411e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=19e-6
mMainBias14 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=13e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=13e-6
mSimpleFirstStageLoad17 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=69e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=284e-6
mSimpleFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=69e-6
mMainBias20 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=23e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_37_9

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 5.13201 mW
** Area: 5401 (mu_m)^2
** Transit frequency: 4.30701 MHz
** Transit frequency with error factor: 4.30503 MHz
** Slew rate: 4.11993 V/mu_s
** Phase margin: 68.755°
** CMRR: 98 dB
** negPSRR: 98 dB
** posPSRR: 94 dB
** VoutMax: 4.25 V
** VoutMin: 1.06001 V
** VcmMax: 4.81001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 8.82901e+06 muA
** NormalTransistorNmos: 1.69211e+07 muA
** NormalTransistorPmos: -2.93069e+07 muA
** NormalTransistorPmos: -9.31999e+06 muA
** NormalTransistorPmos: -9.32099e+06 muA
** NormalTransistorPmos: -9.31999e+06 muA
** NormalTransistorPmos: -9.32099e+06 muA
** NormalTransistorNmos: 1.86381e+07 muA
** NormalTransistorNmos: 1.86391e+07 muA
** NormalTransistorNmos: 9.31901e+06 muA
** NormalTransistorNmos: 9.31901e+06 muA
** NormalTransistorNmos: 9.4275e+08 muA
** DiodeTransistorNmos: 9.42749e+08 muA
** NormalTransistorPmos: -9.42749e+08 muA
** DiodeTransistorNmos: 2.93061e+07 muA
** NormalTransistorNmos: 2.93051e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -8.82999e+06 muA
** DiodeTransistorPmos: -1.69219e+07 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.46601  V
** outSourceVoltageBiasXXnXX1: 0.733001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX0: 3.78201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.589001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** out1: 3.83601  V
** sourceTransconductance: 1.94301  V
** inner: 0.733001  V


.END