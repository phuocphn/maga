** Name: two_stage_single_output_op_amp_52_3

.MACRO two_stage_single_output_op_amp_52_3 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=11e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=17e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=61e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=61e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=34e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=376e-6
mFoldedCascodeFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=95e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=56e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=35e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=35e-6
mSecondStage1StageBias15 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=347e-6
mMainBias16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mMainBias17 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSecondStage1StageBias18 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=596e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=56e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.10001e-12
.EOM two_stage_single_output_op_amp_52_3

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 2.45701 mW
** Area: 7154 (mu_m)^2
** Transit frequency: 4.45601 MHz
** Transit frequency with error factor: 4.45573 MHz
** Slew rate: 3.67197 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 4.02001 V
** VoutMin: 0.310001 V
** VcmMax: 5.17001 V
** VcmMin: 0.790001 V


** Expected Currents: 
** NormalTransistorPmos: -2.53459e+07 muA
** NormalTransistorPmos: -2.33189e+07 muA
** NormalTransistorPmos: -2.25759e+07 muA
** NormalTransistorPmos: -3.54849e+07 muA
** NormalTransistorPmos: -2.25759e+07 muA
** NormalTransistorPmos: -3.54849e+07 muA
** DiodeTransistorNmos: 2.25751e+07 muA
** NormalTransistorNmos: 2.25751e+07 muA
** NormalTransistorNmos: 2.25751e+07 muA
** NormalTransistorNmos: 2.58191e+07 muA
** NormalTransistorNmos: 1.29101e+07 muA
** NormalTransistorNmos: 1.29101e+07 muA
** NormalTransistorNmos: 3.51816e+08 muA
** NormalTransistorPmos: -3.51815e+08 muA
** NormalTransistorPmos: -3.51814e+08 muA
** DiodeTransistorNmos: 2.53451e+07 muA
** DiodeTransistorNmos: 2.33181e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.45301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.927001  V
** inputVoltageBiasXXnXX2: 0.636001  V
** out: 2.5  V
** outFirstStage: 0.719001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.355001  V
** out1: 0.560001  V
** sourceGCC1: 4.16701  V
** sourceGCC2: 4.16701  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 4.19801  V


.END