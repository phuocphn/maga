** Name: one_stage_single_output_op_amp95

.MACRO one_stage_single_output_op_amp95 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=18e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=25e-6
mTelescopicFirstStageLoad3 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=73e-6
mTelescopicFirstStageLoad4 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mTelescopicFirstStageLoad6 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=72e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=18e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=18e-6
mTelescopicFirstStageLoad9 out outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=72e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
mTelescopicFirstStageStageBias11 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=211e-6
mTelescopicFirstStageLoad12 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
mTelescopicFirstStageLoad13 out FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=73e-6
mMainBias14 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=57e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp95

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 0.672001 mW
** Area: 2050 (mu_m)^2
** Transit frequency: 3.63001 MHz
** Transit frequency with error factor: 3.62952 MHz
** Slew rate: 5.78845 V/mu_s
** Phase margin: 86.5167°
** CMRR: 151 dB
** VoutMax: 4.06001 V
** VoutMin: 0.460001 V
** VcmMax: 3.75 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 8.41401e+06 muA
** NormalTransistorPmos: -4.74589e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** DiodeTransistorPmos: -3.42849e+07 muA
** DiodeTransistorPmos: -3.42859e+07 muA
** NormalTransistorPmos: -3.42849e+07 muA
** NormalTransistorPmos: -3.42859e+07 muA
** NormalTransistorNmos: 1.16028e+08 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** DiodeTransistorNmos: 4.74581e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.41499e+06 muA


** Expected Voltages: 
** ibias: 0.567001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 4.13001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerOutputLoad2: 3.49301  V
** innerTransistorStack1Load2: 4.21901  V
** innerTransistorStack2Load2: 4.21901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END