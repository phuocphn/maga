** Name: two_stage_single_output_op_amp_197_10

.MACRO two_stage_single_output_op_amp_197_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=2e-6 W=35e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=19e-6
mMainBias4 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=25e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=172e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=56e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=54e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=19e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=7e-6 W=591e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=35e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=54e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=312e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=344e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=463e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=463e-6
mSimpleFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=276e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=401e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=594e-6
mSimpleFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=276e-6
mMainBias22 outVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=163e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.60001e-12
.EOM two_stage_single_output_op_amp_197_10

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 8.91401 mW
** Area: 14808 (mu_m)^2
** Transit frequency: 4.04701 MHz
** Transit frequency with error factor: 4.04405 MHz
** Slew rate: 3.81454 V/mu_s
** Phase margin: 60.1606°
** CMRR: 125 dB
** VoutMax: 4.54001 V
** VoutMin: 0.210001 V
** VcmMax: 4.75 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 1.62454e+08 muA
** NormalTransistorNmos: 1.80508e+08 muA
** NormalTransistorPmos: -1.71061e+08 muA
** DiodeTransistorNmos: 4.61605e+08 muA
** DiodeTransistorNmos: 4.61604e+08 muA
** NormalTransistorNmos: 4.61605e+08 muA
** NormalTransistorNmos: 4.61604e+08 muA
** NormalTransistorPmos: -4.76297e+08 muA
** NormalTransistorPmos: -4.76298e+08 muA
** NormalTransistorPmos: -4.76297e+08 muA
** NormalTransistorPmos: -4.76298e+08 muA
** NormalTransistorNmos: 2.93851e+07 muA
** NormalTransistorNmos: 2.93841e+07 muA
** NormalTransistorNmos: 1.46931e+07 muA
** NormalTransistorNmos: 1.46931e+07 muA
** NormalTransistorNmos: 3.06143e+08 muA
** NormalTransistorPmos: -3.06142e+08 muA
** NormalTransistorPmos: -3.06143e+08 muA
** DiodeTransistorNmos: 1.71062e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.62453e+08 muA
** DiodeTransistorPmos: -1.80507e+08 muA


** Expected Voltages: 
** ibias: 0.613001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.14301  V
** outVoltageBiasXXnXX1: 0.806001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.09501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.12901  V
** innerStageBias: 0.209001  V
** innerTransistorStack1Load2: 4.56001  V
** innerTransistorStack2Load1: 1.12901  V
** innerTransistorStack2Load2: 4.56001  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.41901  V


.END