** Name: two_stage_single_output_op_amp_24_2

.MACRO two_stage_single_output_op_amp_24_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=35e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=24e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=91e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=257e-6
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=60e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=75e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=75e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=133e-6
mSecondStage1Transconductor10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=535e-6
mSimpleFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=60e-6
mMainBias12 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=16e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=113e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=257e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=91e-6
mMainBias16 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=158e-6
mSecondStage1StageBias17 out ibias sourcePmos sourcePmos pmos4 L=5e-6 W=600e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=113e-6
mMainBias19 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=56e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.8001e-12
.EOM two_stage_single_output_op_amp_24_2

** Expected Performance Values: 
** Gain: 105 dB
** Power consumption: 2.21101 mW
** Area: 12529 (mu_m)^2
** Transit frequency: 3.90501 MHz
** Transit frequency with error factor: 3.90283 MHz
** Slew rate: 4.12803 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** negPSRR: 107 dB
** posPSRR: 196 dB
** VoutMax: 4.66001 V
** VoutMin: 0.300001 V
** VcmMax: 3.16001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.05521e+07 muA
** NormalTransistorPmos: -2.35679e+07 muA
** NormalTransistorPmos: -6.60029e+07 muA
** NormalTransistorNmos: 2.85751e+07 muA
** NormalTransistorNmos: 2.85741e+07 muA
** NormalTransistorNmos: 2.85751e+07 muA
** NormalTransistorNmos: 2.85741e+07 muA
** NormalTransistorPmos: -5.71529e+07 muA
** DiodeTransistorPmos: -5.71539e+07 muA
** NormalTransistorPmos: -2.85759e+07 muA
** NormalTransistorPmos: -2.85759e+07 muA
** NormalTransistorNmos: 2.54834e+08 muA
** NormalTransistorNmos: 2.54833e+08 muA
** NormalTransistorPmos: -2.54833e+08 muA
** DiodeTransistorNmos: 2.35671e+07 muA
** DiodeTransistorNmos: 6.60021e+07 muA
** DiodeTransistorPmos: -2.05529e+07 muA
** NormalTransistorPmos: -2.05529e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.09301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.32401  V
** outSourceVoltageBiasXXpXX1: 4.16201  V
** outVoltageBiasXXnXX0: 0.580001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.23201  V
** innerTransconductance: 0.150001  V
** inner: 4.16201  V


.END