** Name: two_stage_single_output_op_amp_189_11

.MACRO two_stage_single_output_op_amp_189_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=31e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=9e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=38e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=478e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=9e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=31e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=9e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=506e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=391e-6
mMainBias12 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=559e-6
mSecondStage1StageBias13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=522e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=2e-6 W=41e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=9e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=442e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=442e-6
mSimpleFirstStageLoad18 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=465e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=293e-6
mSecondStage1Transconductor20 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
mSimpleFirstStageLoad21 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=465e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_189_11

** Expected Performance Values: 
** Gain: 140 dB
** Power consumption: 12.2211 mW
** Area: 12246 (mu_m)^2
** Transit frequency: 3.97501 MHz
** Transit frequency with error factor: 3.97106 MHz
** Slew rate: 3.80206 V/mu_s
** Phase margin: 64.1713°
** CMRR: 129 dB
** VoutMax: 4.25 V
** VoutMin: 0.710001 V
** VcmMax: 4.66001 V
** VcmMin: 1.33001 V


** Expected Currents: 
** NormalTransistorNmos: 3.85829e+08 muA
** NormalTransistorNmos: 5.50097e+08 muA
** NormalTransistorNmos: 4.91776e+08 muA
** NormalTransistorNmos: 4.91777e+08 muA
** DiodeTransistorNmos: 4.91776e+08 muA
** NormalTransistorPmos: -5.00604e+08 muA
** NormalTransistorPmos: -5.00605e+08 muA
** NormalTransistorPmos: -5.00605e+08 muA
** NormalTransistorPmos: -5.00605e+08 muA
** NormalTransistorNmos: 1.76571e+07 muA
** NormalTransistorNmos: 1.76581e+07 muA
** NormalTransistorNmos: 8.82901e+06 muA
** NormalTransistorNmos: 8.82901e+06 muA
** NormalTransistorNmos: 4.97109e+08 muA
** NormalTransistorNmos: 4.97108e+08 muA
** NormalTransistorPmos: -4.97108e+08 muA
** NormalTransistorPmos: -4.97109e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.85828e+08 muA
** DiodeTransistorPmos: -5.50096e+08 muA


** Expected Voltages: 
** ibias: 1.125  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** inputVoltageBiasXXpXX2: 3.93101  V
** out: 2.5  V
** outFirstStage: 3.90101  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.504001  V
** innerTransistorStack1Load2: 4.49501  V
** innerTransistorStack2Load2: 4.49501  V
** out1: 2.09501  V
** sourceTransconductance: 1.94201  V
** innerStageBias: 0.570001  V
** innerTransconductance: 4.46501  V


.END