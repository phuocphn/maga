** Name: two_stage_single_output_op_amp_105_5

.MACRO two_stage_single_output_op_amp_105_5 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=4e-6 W=14e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=14e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=37e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos4 L=2e-6 W=11e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=69e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=523e-6
mMainBias7 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=9e-6 W=220e-6
mTelescopicFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=4e-6 W=14e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=530e-6
mTelescopicFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=14e-6
mMainBias12 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=159e-6
mMainBias13 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=224e-6
mTelescopicFirstStageStageBias14 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=80e-6
mTelescopicFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=9e-6 W=23e-6
mTelescopicFirstStageTransconductor16 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=53e-6
mTelescopicFirstStageTransconductor17 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=53e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=69e-6
mMainBias19 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mSecondStage1StageBias20 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=523e-6
mTelescopicFirstStageLoad21 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=9e-6 W=23e-6
mTelescopicFirstStageStageBias22 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=338e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_105_5

** Expected Performance Values: 
** Gain: 144 dB
** Power consumption: 5.60801 mW
** Area: 14948 (mu_m)^2
** Transit frequency: 2.68501 MHz
** Transit frequency with error factor: 2.68489 MHz
** Slew rate: 32.5197 V/mu_s
** Phase margin: 60.1606°
** CMRR: 127 dB
** VoutMax: 3 V
** VoutMin: 0.300001 V
** VcmMax: 3 V
** VcmMin: 0.930001 V


** Expected Currents: 
** NormalTransistorNmos: 1.04893e+08 muA
** NormalTransistorNmos: 1.48034e+08 muA
** NormalTransistorPmos: -2.41989e+07 muA
** NormalTransistorPmos: -6.66799e+06 muA
** NormalTransistorPmos: -6.66799e+06 muA
** DiodeTransistorNmos: 6.66701e+06 muA
** DiodeTransistorNmos: 6.66701e+06 muA
** NormalTransistorNmos: 6.66701e+06 muA
** NormalTransistorNmos: 6.66701e+06 muA
** NormalTransistorPmos: -1.61372e+08 muA
** NormalTransistorPmos: -1.61373e+08 muA
** NormalTransistorPmos: -6.66899e+06 muA
** NormalTransistorPmos: -6.66899e+06 muA
** NormalTransistorNmos: 8.11126e+08 muA
** NormalTransistorPmos: -8.11125e+08 muA
** DiodeTransistorPmos: -8.11125e+08 muA
** DiodeTransistorNmos: 2.41981e+07 muA
** DiodeTransistorPmos: -1.04892e+08 muA
** NormalTransistorPmos: -1.04893e+08 muA
** DiodeTransistorPmos: -1.48033e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.07701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.558001  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outInputVoltageBiasXXpXX1: 2.43601  V
** outSourceVoltageBiasXXpXX1: 3.71801  V
** outSourceVoltageBiasXXpXX3: 3.96101  V
** outVoltageBiasXXpXX2: 2.08201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.23101  V
** innerStageBias: 3.87101  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 3.02701  V
** sourceGCC2: 3.02701  V
** inner: 3.71101  V


.END