** Name: one_stage_single_output_op_amp75

.MACRO one_stage_single_output_op_amp75 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=50e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=40e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=17e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=141e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=50e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=85e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=85e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=113e-6
mFoldedCascodeFirstStageLoad11 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=184e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=95e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=111e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=111e-6
mFoldedCascodeFirstStageLoad15 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=95e-6
mMainBias16 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mMainBias17 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp75

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 1.55401 mW
** Area: 5296 (mu_m)^2
** Transit frequency: 3.36501 MHz
** Transit frequency with error factor: 3.36477 MHz
** Slew rate: 3.73915 V/mu_s
** Phase margin: 89.3815°
** CMRR: 139 dB
** VoutMax: 3.99001 V
** VoutMin: 0.470001 V
** VcmMax: 5.17001 V
** VcmMin: 1.43001 V


** Expected Currents: 
** NormalTransistorPmos: -4.43809e+07 muA
** NormalTransistorPmos: -2.12909e+07 muA
** NormalTransistorPmos: -7.50269e+07 muA
** NormalTransistorPmos: -1.12538e+08 muA
** NormalTransistorPmos: -7.50279e+07 muA
** NormalTransistorPmos: -1.12539e+08 muA
** DiodeTransistorNmos: 7.50261e+07 muA
** NormalTransistorNmos: 7.50271e+07 muA
** NormalTransistorNmos: 7.50261e+07 muA
** NormalTransistorNmos: 7.50251e+07 muA
** NormalTransistorNmos: 7.50241e+07 muA
** NormalTransistorNmos: 3.75131e+07 muA
** NormalTransistorNmos: 3.75131e+07 muA
** DiodeTransistorNmos: 4.43801e+07 muA
** DiodeTransistorNmos: 2.12901e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.45301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.07201  V
** outVoltageBiasXXnXX2: 0.629001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.449001  V
** innerTransistorStack2Load2: 0.497001  V
** out1: 0.702001  V
** sourceGCC1: 4.22701  V
** sourceGCC2: 4.22701  V
** sourceTransconductance: 1.91801  V


.END