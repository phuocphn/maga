** Name: two_stage_single_output_op_amp_152_8

.MACRO two_stage_single_output_op_amp_152_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=8e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=110e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=13e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=63e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=548e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=156e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=10e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=63e-6
mSimpleFirstStageLoad14 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=7e-6 W=285e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=65e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=65e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=214e-6
mSimpleFirstStageLoad18 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=285e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=58e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=31e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.90001e-12
.EOM two_stage_single_output_op_amp_152_8

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 6.38401 mW
** Area: 9644 (mu_m)^2
** Transit frequency: 4.23701 MHz
** Transit frequency with error factor: 4.23533 MHz
** Slew rate: 3.99348 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** VoutMax: 4.25 V
** VoutMin: 0.730001 V
** VcmMax: 4.59001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorPmos: -4.54059e+07 muA
** NormalTransistorPmos: -2.37889e+07 muA
** DiodeTransistorNmos: 3.85991e+07 muA
** NormalTransistorNmos: 3.86001e+07 muA
** NormalTransistorNmos: 3.86011e+07 muA
** DiodeTransistorNmos: 3.86001e+07 muA
** NormalTransistorPmos: -5.05999e+07 muA
** NormalTransistorPmos: -5.06009e+07 muA
** NormalTransistorPmos: -5.06019e+07 muA
** NormalTransistorPmos: -5.06009e+07 muA
** NormalTransistorNmos: 2.39991e+07 muA
** NormalTransistorNmos: 1.20001e+07 muA
** NormalTransistorNmos: 1.20001e+07 muA
** NormalTransistorNmos: 1.08642e+09 muA
** NormalTransistorNmos: 1.08642e+09 muA
** NormalTransistorPmos: -1.08641e+09 muA
** DiodeTransistorNmos: 4.54051e+07 muA
** DiodeTransistorNmos: 2.37881e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 3.88501  V
** outVoltageBiasXXnXX1: 1.13401  V
** outVoltageBiasXXnXX2: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerTransistorStack1Load1: 1.08401  V
** innerTransistorStack1Load2: 3.95901  V
** innerTransistorStack2Load1: 1.08301  V
** innerTransistorStack2Load2: 3.95901  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.153001  V


.END