** Name: one_stage_single_output_op_amp60

.MACRO one_stage_single_output_op_amp60 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=5e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=77e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=572e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=51e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=109e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=109e-6
mFoldedCascodeFirstStageLoad9 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=51e-6
mFoldedCascodeFirstStageLoad10 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=185e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=185e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=572e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=77e-6
mMainBias15 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=45e-6
mFoldedCascodeFirstStageLoad16 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp60

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 1.20701 mW
** Area: 8000 (mu_m)^2
** Transit frequency: 2.51201 MHz
** Transit frequency with error factor: 2.51226 MHz
** Slew rate: 3.50002 V/mu_s
** Phase margin: 89.3815°
** CMRR: 126 dB
** VoutMax: 3.53001 V
** VoutMin: 0.740001 V
** VcmMax: 3.29001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -5.88599e+06 muA
** NormalTransistorNmos: 7.00511e+07 muA
** NormalTransistorNmos: 1.0779e+08 muA
** NormalTransistorNmos: 7.00481e+07 muA
** NormalTransistorNmos: 1.07787e+08 muA
** NormalTransistorPmos: -7.00499e+07 muA
** NormalTransistorPmos: -7.00489e+07 muA
** DiodeTransistorPmos: -7.00499e+07 muA
** NormalTransistorPmos: -7.54779e+07 muA
** DiodeTransistorPmos: -7.54769e+07 muA
** NormalTransistorPmos: -3.77389e+07 muA
** NormalTransistorPmos: -3.77389e+07 muA
** DiodeTransistorNmos: 5.88501e+06 muA
** DiodeTransistorNmos: 5.88601e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.52901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.12901  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.26501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.16301  V
** out1: 2.97001  V
** sourceGCC1: 0.543001  V
** sourceGCC2: 0.543001  V
** sourceTransconductance: 3.30201  V
** inner: 4.26301  V


.END