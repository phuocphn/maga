** Name: symmetrical_op_amp115

.MACRO symmetrical_op_amp115 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=17e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=1e-6 W=16e-6
mMainBias4 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=42e-6
mSecondStage1StageBias6 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mSymmetricalFirstStageTransconductor7 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=8e-6
mSecondStage1StageBias8 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=17e-6
mSymmetricalFirstStageTransconductor9 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=8e-6
mMainBias10 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=5e-6 W=169e-6
mSymmetricalFirstStageLoad11 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=17e-6
mSymmetricalFirstStageLoad12 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=17e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=52e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=52e-6
mSymmetricalFirstStageLoad15 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=30e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=93e-6
mSecondStage1Transconductor17 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=93e-6
mSymmetricalFirstStageLoad18 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=30e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp115

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 1.04501 mW
** Area: 2741 (mu_m)^2
** Transit frequency: 2.54901 MHz
** Transit frequency with error factor: 2.54943 MHz
** Slew rate: 3.75003 V/mu_s
** Phase margin: 75.0575°
** CMRR: 141 dB
** negPSRR: 114 dB
** posPSRR: 61 dB
** VoutMax: 4.25 V
** VoutMin: 0.770001 V
** VcmMax: 4.81001 V
** VcmMin: 0.820001 V


** Expected Currents: 
** NormalTransistorNmos: 9.96491e+07 muA
** NormalTransistorPmos: -1.21789e+07 muA
** NormalTransistorPmos: -1.21799e+07 muA
** NormalTransistorPmos: -1.21789e+07 muA
** NormalTransistorPmos: -1.21799e+07 muA
** NormalTransistorNmos: 2.43571e+07 muA
** NormalTransistorNmos: 1.21781e+07 muA
** NormalTransistorNmos: 1.21781e+07 muA
** NormalTransistorNmos: 3.75451e+07 muA
** NormalTransistorNmos: 3.75441e+07 muA
** NormalTransistorPmos: -3.75459e+07 muA
** NormalTransistorPmos: -3.75449e+07 muA
** DiodeTransistorNmos: 3.75431e+07 muA
** DiodeTransistorNmos: 3.75421e+07 muA
** NormalTransistorPmos: -3.75439e+07 muA
** NormalTransistorPmos: -3.75449e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.96499e+07 muA


** Expected Voltages: 
** ibias: 0.591001  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 0.605001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 1.17601  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.86201  V
** innerStageBias: 0.609001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END