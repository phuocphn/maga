** Name: two_stage_single_output_op_amp_79_9

.MACRO two_stage_single_output_op_amp_79_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=56e-6
mSecondStage1StageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=300e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mMainBias4 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=285e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=10e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=24e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=131e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=174e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=174e-6
mFoldedCascodeFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=101e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=58e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=58e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=81e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=56e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=300e-6
mFoldedCascodeFirstStageLoad16 outFirstStage outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=101e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=164e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=119e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=119e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=207e-6
mFoldedCascodeFirstStageLoad21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=164e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=467e-6
mMainBias23 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=81e-6
mMainBias24 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=177e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.80001e-12
.EOM two_stage_single_output_op_amp_79_9

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 7.39501 mW
** Area: 14206 (mu_m)^2
** Transit frequency: 4.49701 MHz
** Transit frequency with error factor: 4.4966 MHz
** Slew rate: 4.84709 V/mu_s
** Phase margin: 60.1606°
** CMRR: 147 dB
** VoutMax: 4.25 V
** VoutMin: 0.810001 V
** VcmMax: 5.19001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorPmos: -1.97321e+08 muA
** NormalTransistorPmos: -3.44239e+07 muA
** NormalTransistorPmos: -7.52229e+07 muA
** NormalTransistorPmos: -3.33029e+07 muA
** NormalTransistorPmos: -5.05729e+07 muA
** NormalTransistorPmos: -3.33029e+07 muA
** NormalTransistorPmos: -5.05729e+07 muA
** NormalTransistorNmos: 3.33021e+07 muA
** NormalTransistorNmos: 3.33011e+07 muA
** NormalTransistorNmos: 3.33021e+07 muA
** NormalTransistorNmos: 3.33011e+07 muA
** NormalTransistorNmos: 3.45371e+07 muA
** NormalTransistorNmos: 3.45361e+07 muA
** NormalTransistorNmos: 1.72691e+07 muA
** NormalTransistorNmos: 1.72691e+07 muA
** NormalTransistorNmos: 1.05088e+09 muA
** DiodeTransistorNmos: 1.05088e+09 muA
** NormalTransistorPmos: -1.05087e+09 muA
** DiodeTransistorNmos: 1.97322e+08 muA
** NormalTransistorNmos: 1.97321e+08 muA
** DiodeTransistorNmos: 3.44231e+07 muA
** DiodeTransistorNmos: 7.52221e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.21601  V
** outSourceVoltageBiasXXnXX1: 0.608001  V
** outSourceVoltageBiasXXpXX1: 4.21901  V
** outVoltageBiasXXnXX2: 0.955001  V
** outVoltageBiasXXnXX3: 0.581001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.376001  V
** innerTransistorStack1Load2: 0.397001  V
** innerTransistorStack2Load2: 0.397001  V
** out1: 0.555001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.91701  V
** inner: 0.606001  V


.END