** Name: two_stage_single_output_op_amp_68_10

.MACRO two_stage_single_output_op_amp_68_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=33e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=9e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=238e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=238e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=57e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=421e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=115e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=66e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=43e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=43e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=289e-6
mFoldedCascodeFirstStageLoad12 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=66e-6
mMainBias13 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=559e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=238e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=24e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=24e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=421e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=507e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=57e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=389e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=238e-6
mMainBias23 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=254e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.20001e-12
.EOM two_stage_single_output_op_amp_68_10

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 10.3851 mW
** Area: 14550 (mu_m)^2
** Transit frequency: 3.91501 MHz
** Transit frequency with error factor: 3.91497 MHz
** Slew rate: 7.19621 V/mu_s
** Phase margin: 60.1606°
** CMRR: 135 dB
** VoutMax: 4.25 V
** VoutMin: 0.160001 V
** VcmMax: 3.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.16765e+09 muA
** NormalTransistorPmos: -4.43589e+07 muA
** NormalTransistorPmos: -6.81759e+07 muA
** NormalTransistorNmos: 5.24341e+07 muA
** NormalTransistorNmos: 8.98881e+07 muA
** NormalTransistorNmos: 5.24301e+07 muA
** NormalTransistorNmos: 8.98821e+07 muA
** DiodeTransistorPmos: -5.24329e+07 muA
** NormalTransistorPmos: -5.24319e+07 muA
** NormalTransistorPmos: -5.24309e+07 muA
** DiodeTransistorPmos: -5.24319e+07 muA
** NormalTransistorPmos: -7.49049e+07 muA
** DiodeTransistorPmos: -7.49039e+07 muA
** NormalTransistorPmos: -3.74529e+07 muA
** NormalTransistorPmos: -3.74529e+07 muA
** NormalTransistorNmos: 5.97041e+08 muA
** NormalTransistorPmos: -5.9704e+08 muA
** NormalTransistorPmos: -5.97041e+08 muA
** DiodeTransistorNmos: 4.43581e+07 muA
** DiodeTransistorNmos: 6.81751e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.16764e+09 muA


** Expected Voltages: 
** ibias: 3.42601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.562001  V
** out: 2.5  V
** outFirstStage: 3.92101  V
** outSourceVoltageBiasXXpXX1: 4.21401  V
** outVoltageBiasXXnXX1: 0.999001  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.27901  V
** innerTransistorStack2Load2: 4.27901  V
** out1: 3.55801  V
** sourceGCC1: 0.357001  V
** sourceGCC2: 0.357001  V
** sourceTransconductance: 3.48001  V
** innerTransconductance: 4.48501  V
** inner: 4.21101  V


.END