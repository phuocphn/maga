** Name: two_stage_single_output_op_amp_76_10

.MACRO two_stage_single_output_op_amp_76_10 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=102e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=36e-6
mMainBias3 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=5e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=89e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=55e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=102e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=34e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=34e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=89e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSecondStage1StageBias13 out inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=244e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=187e-6
mMainBias15 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=321e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=534e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=534e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=400e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=506e-6
mMainBias21 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=192e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=321e-6
mMainBias24 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.8001e-12
.EOM two_stage_single_output_op_amp_76_10

** Expected Performance Values: 
** Gain: 135 dB
** Power consumption: 6.25801 mW
** Area: 14979 (mu_m)^2
** Transit frequency: 4.31201 MHz
** Transit frequency with error factor: 4.31165 MHz
** Slew rate: 4.06362 V/mu_s
** Phase margin: 60.1606°
** CMRR: 149 dB
** VoutMax: 4.25 V
** VoutMin: 0.650001 V
** VcmMax: 5.23001 V
** VcmMin: 1.37001 V


** Expected Currents: 
** NormalTransistorNmos: 3.55351e+07 muA
** NormalTransistorPmos: -3.66499e+06 muA
** NormalTransistorPmos: -9.19379e+07 muA
** NormalTransistorPmos: -3.53779e+07 muA
** NormalTransistorPmos: -6.47589e+07 muA
** NormalTransistorPmos: -9.71369e+07 muA
** NormalTransistorPmos: -6.47619e+07 muA
** NormalTransistorPmos: -9.71419e+07 muA
** DiodeTransistorNmos: 6.47601e+07 muA
** NormalTransistorNmos: 6.47611e+07 muA
** NormalTransistorNmos: 6.47601e+07 muA
** NormalTransistorNmos: 6.47571e+07 muA
** DiodeTransistorNmos: 6.47561e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 8.70761e+08 muA
** NormalTransistorPmos: -8.7076e+08 muA
** NormalTransistorPmos: -8.70761e+08 muA
** DiodeTransistorNmos: 3.66401e+06 muA
** NormalTransistorNmos: 3.66301e+06 muA
** DiodeTransistorNmos: 9.19371e+07 muA
** DiodeTransistorNmos: 3.53771e+07 muA
** DiodeTransistorPmos: -3.55359e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.957001  V
** inputVoltageBiasXXnXX3: 1.05201  V
** out: 2.5  V
** outFirstStage: 4.08701  V
** outInputVoltageBiasXXnXX1: 1.22401  V
** outSourceVoltageBiasXXnXX1: 0.612001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.65101  V
** inner: 0.610001  V


.END