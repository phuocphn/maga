** Name: one_stage_single_output_op_amp51

.MACRO one_stage_single_output_op_amp51 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=66e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=83e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=66e-6
mFoldedCascodeFirstStageTransconductor6 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=39e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=39e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=85e-6
mMainBias9 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=56e-6
mFoldedCascodeFirstStageLoad10 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=47e-6
mFoldedCascodeFirstStageLoad11 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=230e-6
mFoldedCascodeFirstStageLoad12 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=177e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=177e-6
mFoldedCascodeFirstStageLoad14 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=230e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp51

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 1.85101 mW
** Area: 1906 (mu_m)^2
** Transit frequency: 2.94101 MHz
** Transit frequency with error factor: 2.94143 MHz
** Slew rate: 4.65499 V/mu_s
** Phase margin: 88.8085°
** CMRR: 143 dB
** VoutMax: 4.07001 V
** VoutMin: 0.740001 V
** VcmMax: 5.19001 V
** VcmMin: 0.860001 V


** Expected Currents: 
** NormalTransistorNmos: 6.92531e+07 muA
** NormalTransistorPmos: -9.34109e+07 muA
** NormalTransistorPmos: -1.45489e+08 muA
** NormalTransistorPmos: -9.34109e+07 muA
** NormalTransistorPmos: -1.45489e+08 muA
** NormalTransistorNmos: 9.34101e+07 muA
** NormalTransistorNmos: 9.34101e+07 muA
** DiodeTransistorNmos: 9.34101e+07 muA
** NormalTransistorNmos: 1.04158e+08 muA
** NormalTransistorNmos: 5.20781e+07 muA
** NormalTransistorNmos: 5.20781e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.92539e+07 muA
** DiodeTransistorPmos: -6.92529e+07 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.22101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.587001  V
** out1: 1.14501  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.81301  V


.END