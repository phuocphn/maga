** Name: two_stage_single_output_op_amp_13_11

.MACRO two_stage_single_output_op_amp_13_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=213e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=4e-6 W=213e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=35e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=279e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=55e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mMainBias10 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=38e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=589e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=279e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=61e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=213e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=390e-6
mSecondStage1Transconductor16 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=596e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=4e-6 W=213e-6
mMainBias18 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=49e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16e-12
.EOM two_stage_single_output_op_amp_13_11

** Expected Performance Values: 
** Gain: 142 dB
** Power consumption: 8.09601 mW
** Area: 14894 (mu_m)^2
** Transit frequency: 7.04001 MHz
** Transit frequency with error factor: 7.03626 MHz
** Slew rate: 6.68326 V/mu_s
** Phase margin: 60.1606°
** CMRR: 106 dB
** negPSRR: 113 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 0.610001 V
** VcmMax: 3.87001 V
** VcmMin: 0.900001 V


** Expected Currents: 
** NormalTransistorNmos: 7.55331e+07 muA
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorPmos: -1.03955e+08 muA
** DiodeTransistorPmos: -5.39169e+07 muA
** NormalTransistorPmos: -5.39179e+07 muA
** NormalTransistorPmos: -5.39169e+07 muA
** DiodeTransistorPmos: -5.39179e+07 muA
** NormalTransistorNmos: 1.07834e+08 muA
** NormalTransistorNmos: 5.39161e+07 muA
** NormalTransistorNmos: 5.39161e+07 muA
** NormalTransistorNmos: 1.20013e+09 muA
** NormalTransistorNmos: 1.20013e+09 muA
** NormalTransistorPmos: -1.20012e+09 muA
** NormalTransistorPmos: -1.20012e+09 muA
** DiodeTransistorNmos: 1.03956e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.55339e+07 muA
** DiodeTransistorPmos: -1.21839e+08 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.94701  V
** out: 2.5  V
** outFirstStage: 4.02001  V
** outVoltageBiasXXnXX1: 1.01501  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.26701  V
** innerTransistorStack1Load1: 4.26501  V
** out1: 3.46401  V
** sourceTransconductance: 1.94401  V
** innerStageBias: 0.342001  V
** innerTransconductance: 4.58401  V


.END