** Name: two_stage_single_output_op_amp_64_7

.MACRO two_stage_single_output_op_amp_64_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=5e-6 W=167e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=148e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=82e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=278e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=43e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=445e-6
mFoldedCascodeFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=43e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=5e-6 W=167e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=101e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=101e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=278e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=82e-6
mMainBias17 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=239e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=165e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=148e-6
mMainBias20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=521e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_64_7

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 9.35701 mW
** Area: 14931 (mu_m)^2
** Transit frequency: 4.66201 MHz
** Transit frequency with error factor: 4.6617 MHz
** Slew rate: 5.30063 V/mu_s
** Phase margin: 72.1927°
** CMRR: 139 dB
** VoutMax: 4.25 V
** VoutMin: 0.300001 V
** VcmMax: 3.21001 V
** VcmMin: -0.269999 V


** Expected Currents: 
** NormalTransistorPmos: -6.38909e+07 muA
** NormalTransistorPmos: -2.95729e+07 muA
** NormalTransistorNmos: 2.41261e+07 muA
** NormalTransistorNmos: 4.13601e+07 muA
** NormalTransistorNmos: 2.41221e+07 muA
** NormalTransistorNmos: 4.13541e+07 muA
** DiodeTransistorPmos: -2.4125e+07 muA
** DiodeTransistorPmos: -2.41239e+07 muA
** NormalTransistorPmos: -2.41229e+07 muA
** NormalTransistorPmos: -2.41239e+07 muA
** NormalTransistorPmos: -3.44649e+07 muA
** DiodeTransistorPmos: -3.44639e+07 muA
** NormalTransistorPmos: -1.72329e+07 muA
** NormalTransistorPmos: -1.72329e+07 muA
** NormalTransistorNmos: 1.67532e+09 muA
** NormalTransistorPmos: -1.67531e+09 muA
** DiodeTransistorNmos: 6.38901e+07 muA
** DiodeTransistorNmos: 2.95721e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.46401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.702001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.23301  V
** outVoltageBiasXXnXX1: 1.06501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.23401  V
** innerTransistorStack2Load2: 4.23301  V
** out1: 3.45601  V
** sourceGCC1: 0.497001  V
** sourceGCC2: 0.497001  V
** sourceTransconductance: 3.32201  V
** inner: 4.23001  V


.END