** Name: two_stage_single_output_op_amp_195_12

.MACRO two_stage_single_output_op_amp_195_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=27e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=49e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=8e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=23e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=310e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mSecondStage1StageBias7 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=155e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=246e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=27e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=124e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=79e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mMainBias14 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=574e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=310e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=49e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=124e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=196e-6
mSimpleFirstStageLoad19 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=526e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=556e-6
mSecondStage1Transconductor21 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=526e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=175e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.5e-12
.EOM two_stage_single_output_op_amp_195_12

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 12.8081 mW
** Area: 9479 (mu_m)^2
** Transit frequency: 6.06001 MHz
** Transit frequency with error factor: 6.04355 MHz
** Slew rate: 5.71148 V/mu_s
** Phase margin: 60.1606°
** CMRR: 94 dB
** VoutMax: 4.25 V
** VoutMin: 0.870001 V
** VcmMax: 5.22001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 2.74142e+08 muA
** NormalTransistorNmos: 9.36951e+07 muA
** NormalTransistorPmos: -1.05785e+08 muA
** DiodeTransistorNmos: 2.54579e+08 muA
** DiodeTransistorNmos: 2.5458e+08 muA
** NormalTransistorNmos: 2.54579e+08 muA
** NormalTransistorNmos: 2.5458e+08 muA
** NormalTransistorPmos: -3.13622e+08 muA
** NormalTransistorPmos: -3.13622e+08 muA
** NormalTransistorNmos: 1.18088e+08 muA
** NormalTransistorNmos: 1.18087e+08 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorNmos: 1.45079e+09 muA
** DiodeTransistorNmos: 1.45079e+09 muA
** NormalTransistorPmos: -1.45078e+09 muA
** NormalTransistorPmos: -1.45078e+09 muA
** DiodeTransistorNmos: 1.05786e+08 muA
** NormalTransistorNmos: 1.05785e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.74141e+08 muA
** DiodeTransistorPmos: -9.36959e+07 muA


** Expected Voltages: 
** ibias: 1.20201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.05201  V
** outInputVoltageBiasXXnXX1: 1.27801  V
** outSourceVoltageBiasXXnXX1: 0.639001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX2: 4.25301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.530001  V
** innerTransistorStack2Load1: 1.15501  V
** out1: 2.11601  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.61601  V
** inner: 0.639001  V


.END