** Name: two_stage_single_output_op_amp_52_4

.MACRO two_stage_single_output_op_amp_52_4 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=165e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=183e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=23e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=165e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=70e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=70e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=169e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=219e-6
mSecondStage1Transconductor11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=477e-6
mFoldedCascodeFirstStageLoad12 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=54e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=156e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=106e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=106e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=460e-6
mSecondStage1StageBias17 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=598e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=156e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=79e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=94e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.1001e-12
.EOM two_stage_single_output_op_amp_52_4

** Expected Performance Values: 
** Gain: 189 dB
** Power consumption: 4.38201 mW
** Area: 7969 (mu_m)^2
** Transit frequency: 6.66501 MHz
** Transit frequency with error factor: 6.66469 MHz
** Slew rate: 4.45431 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 3.99001 V
** VoutMin: 0.310001 V
** VcmMax: 5.17001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorPmos: -7.96819e+07 muA
** NormalTransistorPmos: -9.53039e+07 muA
** NormalTransistorPmos: -6.30299e+07 muA
** NormalTransistorPmos: -1.0747e+08 muA
** NormalTransistorPmos: -6.30299e+07 muA
** NormalTransistorPmos: -1.0747e+08 muA
** DiodeTransistorNmos: 6.30291e+07 muA
** NormalTransistorNmos: 6.30291e+07 muA
** NormalTransistorNmos: 6.30291e+07 muA
** NormalTransistorNmos: 8.88831e+07 muA
** NormalTransistorNmos: 4.44421e+07 muA
** NormalTransistorNmos: 4.44421e+07 muA
** NormalTransistorNmos: 4.66385e+08 muA
** NormalTransistorNmos: 4.66384e+08 muA
** NormalTransistorPmos: -4.66384e+08 muA
** NormalTransistorPmos: -4.66383e+08 muA
** DiodeTransistorNmos: 7.96811e+07 muA
** DiodeTransistorNmos: 9.53031e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.563001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.921001  V
** outVoltageBiasXXnXX2: 0.627001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.19301  V
** sourceGCC2: 4.19301  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 4.25101  V
** innerTransconductance: 0.364001  V


.END