** Name: symmetrical_op_amp69

.MACRO symmetrical_op_amp69 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=30e-6
mSecondStage1StageBias2 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=24e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mSecondStage1StageBias4 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSymmetricalFirstStageLoad5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=55e-6
mSymmetricalFirstStageLoad6 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=55e-6
mSymmetricalFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=600e-6
mSymmetricalFirstStageStageBias8 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=251e-6
mMainBias9 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=37e-6
mSymmetricalFirstStageTransconductor10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=47e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias11 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=24e-6
mSecondStage1StageBias12 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos4 L=6e-6 W=31e-6
mSymmetricalFirstStageTransconductor13 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=47e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=57e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=57e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=4e-6 W=97e-6
mSecondStage1Transconductor17 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=97e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp69

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 1.82001 mW
** Area: 8404 (mu_m)^2
** Transit frequency: 6.71501 MHz
** Transit frequency with error factor: 6.71527 MHz
** Slew rate: 8.82055 V/mu_s
** Phase margin: 77.3494°
** CMRR: 139 dB
** negPSRR: 57 dB
** posPSRR: 47 dB
** VoutMax: 4.26001 V
** VoutMin: 1.40001 V
** VcmMax: 4.55001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01521e+07 muA
** DiodeTransistorPmos: -8.35559e+07 muA
** DiodeTransistorPmos: -8.35559e+07 muA
** NormalTransistorNmos: 1.6711e+08 muA
** NormalTransistorNmos: 1.67109e+08 muA
** NormalTransistorNmos: 8.35551e+07 muA
** NormalTransistorNmos: 8.35551e+07 muA
** NormalTransistorNmos: 8.83281e+07 muA
** DiodeTransistorNmos: 8.83271e+07 muA
** NormalTransistorPmos: -8.83289e+07 muA
** NormalTransistorPmos: -8.83279e+07 muA
** NormalTransistorNmos: 8.83281e+07 muA
** NormalTransistorPmos: -8.83289e+07 muA
** NormalTransistorPmos: -8.83279e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.01529e+07 muA


** Expected Voltages: 
** ibias: 1.12701  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 4.14301  V
** inStageBiasComplementarySecondStage: 0.954001  V
** innerComplementarySecondStage: 1.80701  V
** out: 2.5  V
** outFirstStage: 4.14301  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.487001  V
** sourceTransconductance: 1.89001  V
** innerTransconductance: 4.70001  V
** inner: 4.70001  V


.END