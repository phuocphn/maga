** Name: one_stage_single_output_op_amp44

.MACRO one_stage_single_output_op_amp44 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=6e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=10e-6 W=82e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=103e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=226e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=226e-6
mFoldedCascodeFirstStageLoad8 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=103e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=141e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=141e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=10e-6 W=586e-6
mMainBias13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=10e-6 W=27e-6
mFoldedCascodeFirstStageLoad14 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=85e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp44

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 1.20201 mW
** Area: 10402 (mu_m)^2
** Transit frequency: 3.39601 MHz
** Transit frequency with error factor: 3.39618 MHz
** Slew rate: 3.60574 V/mu_s
** Phase margin: 87.0896°
** CMRR: 139 dB
** VoutMax: 3.64001 V
** VoutMin: 0.740001 V
** VcmMax: 4.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -3.33399e+06 muA
** NormalTransistorNmos: 7.22751e+07 muA
** NormalTransistorNmos: 1.08579e+08 muA
** NormalTransistorNmos: 7.22751e+07 muA
** NormalTransistorNmos: 1.08579e+08 muA
** NormalTransistorPmos: -7.22759e+07 muA
** NormalTransistorPmos: -7.22759e+07 muA
** DiodeTransistorPmos: -7.22759e+07 muA
** NormalTransistorPmos: -7.26079e+07 muA
** NormalTransistorPmos: -3.63039e+07 muA
** NormalTransistorPmos: -3.63039e+07 muA
** DiodeTransistorNmos: 3.33301e+06 muA
** DiodeTransistorNmos: 3.33401e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.12201  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 3.94601  V
** out1: 3.07201  V
** sourceGCC1: 0.534001  V
** sourceGCC2: 0.534001  V
** sourceTransconductance: 3.23301  V


.END