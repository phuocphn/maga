** Name: two_stage_single_output_op_amp_8_8

.MACRO two_stage_single_output_op_amp_8_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=9e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=46e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=19e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=22e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=385e-6
mSecondStage1StageBias8 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=281e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=19e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mMainBias11 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=150e-6
mSecondStage1Transconductor12 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=254e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=9e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.20001e-12
.EOM two_stage_single_output_op_amp_8_8

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 3.77601 mW
** Area: 3574 (mu_m)^2
** Transit frequency: 3.93901 MHz
** Transit frequency with error factor: 3.92865 MHz
** Slew rate: 6.94169 V/mu_s
** Phase margin: 60.1606°
** CMRR: 83 dB
** negPSRR: 128 dB
** posPSRR: 82 dB
** VoutMax: 4.25 V
** VoutMin: 0.430001 V
** VcmMax: 4.09001 V
** VcmMin: 0.880001 V


** Expected Currents: 
** NormalTransistorNmos: 1.50781e+07 muA
** NormalTransistorPmos: -4.92109e+07 muA
** DiodeTransistorPmos: -1.80729e+07 muA
** NormalTransistorPmos: -1.80729e+07 muA
** NormalTransistorNmos: 3.61441e+07 muA
** NormalTransistorNmos: 1.80721e+07 muA
** NormalTransistorNmos: 1.80721e+07 muA
** NormalTransistorNmos: 6.44741e+08 muA
** NormalTransistorNmos: 6.4474e+08 muA
** NormalTransistorPmos: -6.4474e+08 muA
** DiodeTransistorNmos: 4.92101e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.50789e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.843001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 4.16401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.68601  V
** sourceTransconductance: 1.81401  V
** innerStageBias: 0.205001  V


.END