** Name: two_stage_single_output_op_amp_124_8

.MACRO two_stage_single_output_op_amp_124_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=3e-6 W=6e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=35e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=286e-6
mTelescopicFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=296e-6
mMainBias5 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mTelescopicFirstStageLoad6 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=157e-6
mTelescopicFirstStageLoad7 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=157e-6
mMainBias8 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=33e-6
mTelescopicFirstStageLoad9 FirstStageYinnerOutputLoad2 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=20e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=20e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=20e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=3e-6 W=398e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=286e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=3e-6 W=26e-6
mSecondStage1StageBias15 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=418e-6
mTelescopicFirstStageLoad16 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=20e-6
mTelescopicFirstStageStageBias17 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=296e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=157e-6
mMainBias19 inputVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=174e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=303e-6
mTelescopicFirstStageLoad21 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=5e-6 W=157e-6
mMainBias22 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=215e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.5e-12
.EOM two_stage_single_output_op_amp_124_8

** Expected Performance Values: 
** Gain: 149 dB
** Power consumption: 2.57401 mW
** Area: 14924 (mu_m)^2
** Transit frequency: 2.55201 MHz
** Transit frequency with error factor: 2.55218 MHz
** Slew rate: 8.65507 V/mu_s
** Phase margin: 60.1606°
** CMRR: 144 dB
** VoutMax: 4.69001 V
** VoutMin: 0.710001 V
** VcmMax: 3.81001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 1.70211e+07 muA
** NormalTransistorPmos: -1.08945e+08 muA
** NormalTransistorPmos: -8.80039e+07 muA
** NormalTransistorNmos: 1.26981e+07 muA
** NormalTransistorNmos: 1.26981e+07 muA
** DiodeTransistorPmos: -1.26989e+07 muA
** NormalTransistorPmos: -1.26999e+07 muA
** NormalTransistorPmos: -1.26989e+07 muA
** DiodeTransistorPmos: -1.26999e+07 muA
** NormalTransistorNmos: 1.13399e+08 muA
** DiodeTransistorNmos: 1.13398e+08 muA
** NormalTransistorNmos: 1.26981e+07 muA
** NormalTransistorNmos: 1.26981e+07 muA
** NormalTransistorNmos: 2.65379e+08 muA
** NormalTransistorNmos: 2.65378e+08 muA
** NormalTransistorPmos: -2.65378e+08 muA
** DiodeTransistorNmos: 1.08946e+08 muA
** NormalTransistorNmos: 1.08946e+08 muA
** DiodeTransistorNmos: 8.80031e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.70219e+07 muA


** Expected Voltages: 
** ibias: 1.20501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 2.65001  V
** inputVoltageBiasXXpXX0: 4.05801  V
** out: 2.5  V
** outFirstStage: 4.12201  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX3: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerOutputLoad2: 3.55801  V
** innerSourceLoad2: 4.27201  V
** innerTransistorStack1Load2: 4.27201  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.650001  V
** inner: 0.555001  V


.END