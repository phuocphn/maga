** Name: two_stage_single_output_op_amp_33_9

.MACRO two_stage_single_output_op_amp_33_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=8e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=46e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=234e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=14e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=384e-6
mMainBias7 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=48e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=14e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=30e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=14e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=46e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=387e-6
mMainBias13 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=93e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=234e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=14e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=14e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=468e-6
mSimpleFirstStageLoad18 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=8e-6 W=199e-6
mMainBias19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=351e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_33_9

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 8.82801 mW
** Area: 9388 (mu_m)^2
** Transit frequency: 3.80201 MHz
** Transit frequency with error factor: 3.80075 MHz
** Slew rate: 4.39069 V/mu_s
** Phase margin: 74.4846°
** CMRR: 96 dB
** negPSRR: 108 dB
** posPSRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 1.49001 V
** VcmMax: 4.09001 V
** VcmMin: 1.37001 V


** Expected Currents: 
** NormalTransistorNmos: 2.53093e+08 muA
** NormalTransistorNmos: 6.09191e+07 muA
** NormalTransistorPmos: -2.33654e+08 muA
** DiodeTransistorPmos: -1.00089e+07 muA
** NormalTransistorPmos: -1.00089e+07 muA
** NormalTransistorPmos: -1.00089e+07 muA
** NormalTransistorNmos: 2.00151e+07 muA
** NormalTransistorNmos: 2.00141e+07 muA
** NormalTransistorNmos: 1.00081e+07 muA
** NormalTransistorNmos: 1.00081e+07 muA
** NormalTransistorNmos: 1.18795e+09 muA
** DiodeTransistorNmos: 1.18795e+09 muA
** NormalTransistorPmos: -1.18794e+09 muA
** DiodeTransistorNmos: 2.33655e+08 muA
** NormalTransistorNmos: 2.33654e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.53092e+08 muA
** DiodeTransistorPmos: -6.09199e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.24301  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.90001  V
** outSourceVoltageBiasXXnXX1: 0.950001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.83601  V
** innerStageBias: 0.542001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.91101  V
** inner: 0.945001  V


.END