** Name: two_stage_single_output_op_amp_203_10

.MACRO two_stage_single_output_op_amp_203_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=17e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=14e-6
mMainBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=141e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=101e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=53e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=60e-6
mMainBias11 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=132e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=517e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=17e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=53e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=186e-6
mSimpleFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=194e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=484e-6
mMainBias18 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=194e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=486e-6
mSimpleFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=194e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_203_10

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 5.71401 mW
** Area: 8371 (mu_m)^2
** Transit frequency: 4.72301 MHz
** Transit frequency with error factor: 4.68414 MHz
** Slew rate: 4.48367 V/mu_s
** Phase margin: 70.4739°
** CMRR: 95 dB
** VoutMax: 4.59001 V
** VoutMin: 0.160001 V
** VcmMax: 5.01001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 1.31994e+08 muA
** NormalTransistorNmos: 9.48151e+07 muA
** NormalTransistorPmos: -1.82121e+08 muA
** DiodeTransistorNmos: 1.69096e+08 muA
** NormalTransistorNmos: 1.69097e+08 muA
** NormalTransistorNmos: 1.69096e+08 muA
** DiodeTransistorNmos: 1.69097e+08 muA
** NormalTransistorPmos: -1.79336e+08 muA
** NormalTransistorPmos: -1.79336e+08 muA
** NormalTransistorNmos: 2.04821e+07 muA
** NormalTransistorNmos: 2.04831e+07 muA
** NormalTransistorNmos: 1.02411e+07 muA
** NormalTransistorNmos: 1.02411e+07 muA
** NormalTransistorNmos: 3.6515e+08 muA
** NormalTransistorPmos: -3.65149e+08 muA
** NormalTransistorPmos: -3.6515e+08 muA
** DiodeTransistorNmos: 1.82122e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.31993e+08 muA
** DiodeTransistorPmos: -9.48159e+07 muA


** Expected Voltages: 
** ibias: 0.564001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.732001  V
** inputVoltageBiasXXpXX2: 4.04101  V
** out: 2.5  V
** outFirstStage: 4.23001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.09401  V
** innerStageBias: 0.159001  V
** innerTransistorStack1Load1: 1.09401  V
** out1: 2.09501  V
** sourceTransconductance: 1.94401  V
** innerTransconductance: 4.45501  V


.END