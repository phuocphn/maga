** Name: two_stage_single_output_op_amp_168_6

.MACRO two_stage_single_output_op_amp_168_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=116e-6
mSecondStage1StageBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=30e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=235e-6
mMainBias5 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=1e-6 W=23e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=405e-6
mSimpleFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=322e-6
mSecondStage1StageBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=574e-6
mSimpleFirstStageLoad9 FirstStageYout1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=91e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=264e-6
mSecondStage1Transconductor11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=397e-6
mSimpleFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=91e-6
mMainBias13 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=48e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=30e-6
mSimpleFirstStageTransconductor15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=44e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=322e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=405e-6
mMainBias18 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mMainBias19 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=504e-6
mSecondStage1StageBias20 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=574e-6
mSimpleFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=235e-6
mSimpleFirstStageTransconductor22 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=44e-6
mMainBias23 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=402e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18e-12
.EOM two_stage_single_output_op_amp_168_6

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 5.53601 mW
** Area: 11339 (mu_m)^2
** Transit frequency: 2.95801 MHz
** Transit frequency with error factor: 2.94865 MHz
** Slew rate: 3.97311 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.12001 V
** VoutMin: 0.300001 V
** VcmMax: 3.21001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 9.14231e+07 muA
** NormalTransistorPmos: -1.76005e+08 muA
** NormalTransistorPmos: -2.20937e+08 muA
** DiodeTransistorPmos: -1.37398e+08 muA
** DiodeTransistorPmos: -1.37399e+08 muA
** NormalTransistorPmos: -1.37398e+08 muA
** NormalTransistorPmos: -1.37399e+08 muA
** NormalTransistorNmos: 1.73322e+08 muA
** NormalTransistorNmos: 1.73322e+08 muA
** NormalTransistorPmos: -7.18469e+07 muA
** DiodeTransistorPmos: -7.18479e+07 muA
** NormalTransistorPmos: -3.59229e+07 muA
** NormalTransistorPmos: -3.59229e+07 muA
** NormalTransistorNmos: 2.52148e+08 muA
** NormalTransistorNmos: 2.52147e+08 muA
** NormalTransistorPmos: -2.52145e+08 muA
** DiodeTransistorPmos: -2.52144e+08 muA
** DiodeTransistorNmos: 1.76006e+08 muA
** DiodeTransistorNmos: 2.20938e+08 muA
** DiodeTransistorPmos: -9.14239e+07 muA
** NormalTransistorPmos: -9.14249e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.55901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.42401  V
** outSourceVoltageBiasXXpXX1: 4.21201  V
** outSourceVoltageBiasXXpXX2: 4.28001  V
** outVoltageBiasXXnXX1: 0.705001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.71701  V
** innerTransistorStack2Load1: 3.71501  V
** out1: 2.89601  V
** sourceTransconductance: 3.27701  V
** innerTransconductance: 0.150001  V
** inner: 4.21201  V
** inner: 4.27901  V


.END