** Name: two_stage_single_output_op_amp_203_9

.MACRO two_stage_single_output_op_amp_203_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=9e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=4e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=6e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=511e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mMainBias7 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=101e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=50e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=60e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=511e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=2e-6 W=9e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=50e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=308e-6
mMainBias17 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=264e-6
mSimpleFirstStageLoad19 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=308e-6
mMainBias20 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=61e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.80001e-12
.EOM two_stage_single_output_op_amp_203_9

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 14.9931 mW
** Area: 3881 (mu_m)^2
** Transit frequency: 11.3691 MHz
** Transit frequency with error factor: 11.3391 MHz
** Slew rate: 10.7149 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 1.10001 V
** VcmMax: 5.24001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorPmos: -3.04749e+07 muA
** NormalTransistorPmos: -9.54599e+06 muA
** DiodeTransistorNmos: 1.0795e+08 muA
** NormalTransistorNmos: 1.07951e+08 muA
** NormalTransistorNmos: 1.07952e+08 muA
** DiodeTransistorNmos: 1.07951e+08 muA
** NormalTransistorPmos: -1.55565e+08 muA
** NormalTransistorPmos: -1.55565e+08 muA
** NormalTransistorNmos: 9.52311e+07 muA
** NormalTransistorNmos: 9.52301e+07 muA
** NormalTransistorNmos: 4.76161e+07 muA
** NormalTransistorNmos: 4.76161e+07 muA
** NormalTransistorNmos: 2.62747e+09 muA
** DiodeTransistorNmos: 2.62747e+09 muA
** NormalTransistorPmos: -2.62746e+09 muA
** DiodeTransistorNmos: 3.04741e+07 muA
** NormalTransistorNmos: 3.04731e+07 muA
** DiodeTransistorNmos: 9.54501e+06 muA
** DiodeTransistorNmos: 9.54401e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.28301  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.50401  V
** outSourceVoltageBiasXXnXX1: 0.752001  V
** outSourceVoltageBiasXXnXX2: 0.588001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.640001  V
** innerTransistorStack1Load1: 1.15601  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 0.751001  V


.END