** Name: two_stage_single_output_op_amp_48_7

.MACRO two_stage_single_output_op_amp_48_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=598e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=225e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=186e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=186e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=599e-6
mFoldedCascodeFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=225e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=27e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=27e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=497e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mMainBias16 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=33e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=342e-6
mFoldedCascodeFirstStageLoad18 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=598e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14e-12
.EOM two_stage_single_output_op_amp_48_7

** Expected Performance Values: 
** Gain: 111 dB
** Power consumption: 14.9991 mW
** Area: 6165 (mu_m)^2
** Transit frequency: 7.43901 MHz
** Transit frequency with error factor: 7.43831 MHz
** Slew rate: 22.7068 V/mu_s
** Phase margin: 60.1606°
** CMRR: 129 dB
** VoutMax: 4.45001 V
** VoutMin: 0.190001 V
** VcmMax: 3.52001 V
** VcmMin: -0.379999 V


** Expected Currents: 
** NormalTransistorPmos: -3.55209e+07 muA
** NormalTransistorPmos: -2.98219e+07 muA
** NormalTransistorNmos: 3.23058e+08 muA
** NormalTransistorNmos: 5.52161e+08 muA
** NormalTransistorNmos: 3.23059e+08 muA
** NormalTransistorNmos: 5.52162e+08 muA
** DiodeTransistorPmos: -3.23057e+08 muA
** NormalTransistorPmos: -3.23058e+08 muA
** NormalTransistorPmos: -3.23058e+08 muA
** DiodeTransistorPmos: -3.23058e+08 muA
** NormalTransistorPmos: -4.58206e+08 muA
** NormalTransistorPmos: -2.29103e+08 muA
** NormalTransistorPmos: -2.29103e+08 muA
** NormalTransistorNmos: 1.81024e+09 muA
** NormalTransistorPmos: -1.81023e+09 muA
** DiodeTransistorNmos: 3.55201e+07 muA
** DiodeTransistorNmos: 2.98211e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.05301  V
** inputVoltageBiasXXnXX2: 0.593001  V
** out: 2.5  V
** outFirstStage: 3.89001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.26301  V
** innerTransistorStack1Load2: 4.26301  V
** out1: 3.52601  V
** sourceGCC1: 0.388001  V
** sourceGCC2: 0.388001  V
** sourceTransconductance: 3.75  V


.END