** Name: two_stage_single_output_op_amp_177_6

.MACRO two_stage_single_output_op_amp_177_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=12e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=8e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=469e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad9 FirstStageYinnerOutputLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=201e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=378e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=378e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mSecondStage1Transconductor13 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad14 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=201e-6
mMainBias15 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mSimpleFirstStageTransconductor16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=537e-6
mSimpleFirstStageStageBias17 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mSimpleFirstStageStageBias19 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=330e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=469e-6
mSimpleFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=12e-6
mSimpleFirstStageTransconductor23 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=537e-6
mMainBias24 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=164e-6
mMainBias25 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.3001e-12
.EOM two_stage_single_output_op_amp_177_6

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 14.9831 mW
** Area: 9505 (mu_m)^2
** Transit frequency: 16.1151 MHz
** Transit frequency with error factor: 16.1002 MHz
** Slew rate: 31.2228 V/mu_s
** Phase margin: 60.1606°
** CMRR: 78 dB
** VoutMax: 3.08001 V
** VoutMin: 0.390001 V
** VcmMax: 3.01001 V
** VcmMin: -0.239999 V


** Expected Currents: 
** NormalTransistorNmos: 3.26271e+07 muA
** NormalTransistorPmos: -1.66275e+08 muA
** NormalTransistorPmos: -1.00219e+07 muA
** DiodeTransistorPmos: -1.21839e+08 muA
** NormalTransistorPmos: -1.21839e+08 muA
** NormalTransistorPmos: -1.21839e+08 muA
** DiodeTransistorPmos: -1.21839e+08 muA
** NormalTransistorNmos: 4.26004e+08 muA
** NormalTransistorNmos: 4.26003e+08 muA
** NormalTransistorNmos: 4.26004e+08 muA
** NormalTransistorNmos: 4.26003e+08 muA
** NormalTransistorPmos: -6.08327e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorNmos: 1.91562e+09 muA
** NormalTransistorNmos: 1.91562e+09 muA
** NormalTransistorPmos: -1.91561e+09 muA
** DiodeTransistorPmos: -1.91561e+09 muA
** DiodeTransistorNmos: 1.66276e+08 muA
** DiodeTransistorNmos: 1.00211e+07 muA
** DiodeTransistorPmos: -3.26279e+07 muA
** NormalTransistorPmos: -3.26289e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.599001  V
** outInputVoltageBiasXXpXX1: 2.51401  V
** outSourceVoltageBiasXXpXX1: 3.75701  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX1: 0.793001  V
** outVoltageBiasXXnXX2: 0.568001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerSourceLoad1: 3.68601  V
** innerStageBias: 4.28201  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.229001  V
** innerTransistorStack2Load2: 0.229001  V
** sourceTransconductance: 3.37101  V
** innerTransconductance: 0.194001  V
** inner: 3.75101  V


.END