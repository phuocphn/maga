** Name: two_stage_single_output_op_amp_68_4

.MACRO two_stage_single_output_op_amp_68_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=242e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=6e-6 W=43e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=6e-6 W=95e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=18e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=127e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=147e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=147e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=389e-6
mSecondStage1Transconductor13 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=26e-6
mFoldedCascodeFirstStageLoad14 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=14e-6
mMainBias15 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=14e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=39e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=39e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=127e-6
mSecondStage1StageBias20 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=55e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=18e-6
mMainBias22 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=39e-6
mSecondStage1StageBias23 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=6e-6 W=597e-6
mFoldedCascodeFirstStageLoad24 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=43e-6
mMainBias25 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=151e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_68_4

** Expected Performance Values: 
** Gain: 177 dB
** Power consumption: 2.59201 mW
** Area: 14704 (mu_m)^2
** Transit frequency: 2.57001 MHz
** Transit frequency with error factor: 2.56952 MHz
** Slew rate: 3.77568 V/mu_s
** Phase margin: 62.4525°
** CMRR: 128 dB
** VoutMax: 3.46001 V
** VoutMin: 0.360001 V
** VcmMax: 3.13001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.81001e+06 muA
** NormalTransistorPmos: -2.55526e+08 muA
** NormalTransistorPmos: -6.59969e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 3.99981e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 3.99981e+07 muA
** DiodeTransistorPmos: -2.66659e+07 muA
** NormalTransistorPmos: -2.66669e+07 muA
** NormalTransistorPmos: -2.66659e+07 muA
** DiodeTransistorPmos: -2.66669e+07 muA
** NormalTransistorPmos: -2.66689e+07 muA
** DiodeTransistorPmos: -2.66699e+07 muA
** NormalTransistorPmos: -1.33339e+07 muA
** NormalTransistorPmos: -1.33339e+07 muA
** NormalTransistorNmos: 9.30721e+07 muA
** NormalTransistorNmos: 9.30711e+07 muA
** NormalTransistorPmos: -9.30729e+07 muA
** NormalTransistorPmos: -9.30719e+07 muA
** DiodeTransistorNmos: 2.55527e+08 muA
** DiodeTransistorNmos: 6.59961e+07 muA
** DiodeTransistorPmos: -3.81099e+06 muA
** NormalTransistorPmos: -3.81199e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.93401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.49601  V
** outSourceVoltageBiasXXpXX1: 4.24801  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX1: 0.905001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.24601  V
** innerTransistorStack2Load2: 4.24901  V
** out1: 3.22701  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.42901  V
** innerStageBias: 3.72601  V
** innerTransconductance: 0.294001  V
** inner: 4.24801  V


.END