** Name: symmetrical_op_amp144

.MACRO symmetrical_op_amp144 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=82e-6
mMainBias4 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mSymmetricalFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=80e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=80e-6
mMainBias9 inOutputStageBiasComplementarySecondStage outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=93e-6
mSymmetricalFirstStageLoad10 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=116e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=194e-6
mSecondStage1Transconductor12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=194e-6
mSymmetricalFirstStageLoad13 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=116e-6
mSymmetricalFirstStageStageBias14 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=600e-6
mSymmetricalFirstStageStageBias15 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=185e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=124e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias17 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=124e-6
mSymmetricalFirstStageTransconductor18 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=87e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias19 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=1e-6 W=189e-6
mSecondStage1StageBias20 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=74e-6
mSymmetricalFirstStageTransconductor21 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=87e-6
mMainBias22 out2FirstStage ibias sourcePmos sourcePmos pmos4 L=6e-6 W=115e-6
mMainBias23 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=233e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp144

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 2.31001 mW
** Area: 11953 (mu_m)^2
** Transit frequency: 7.82701 MHz
** Transit frequency with error factor: 7.82727 MHz
** Slew rate: 7.59605 V/mu_s
** Phase margin: 68.755°
** CMRR: 152 dB
** negPSRR: 54 dB
** posPSRR: 72 dB
** VoutMax: 4.58001 V
** VoutMin: 0.320001 V
** VcmMax: 3.37001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.72607e+08 muA
** NormalTransistorPmos: -2.83229e+07 muA
** NormalTransistorPmos: -1.42559e+07 muA
** NormalTransistorNmos: 3.71921e+07 muA
** NormalTransistorNmos: 3.71911e+07 muA
** NormalTransistorNmos: 3.71921e+07 muA
** NormalTransistorNmos: 3.71911e+07 muA
** NormalTransistorPmos: -7.43849e+07 muA
** NormalTransistorPmos: -7.43839e+07 muA
** NormalTransistorPmos: -3.71929e+07 muA
** NormalTransistorPmos: -3.71929e+07 muA
** NormalTransistorNmos: 7.61851e+07 muA
** NormalTransistorNmos: 7.61861e+07 muA
** NormalTransistorPmos: -7.61859e+07 muA
** NormalTransistorPmos: -7.61869e+07 muA
** NormalTransistorPmos: -7.61859e+07 muA
** NormalTransistorPmos: -7.61869e+07 muA
** NormalTransistorNmos: 7.61851e+07 muA
** NormalTransistorNmos: 7.61861e+07 muA
** DiodeTransistorNmos: 2.83221e+07 muA
** DiodeTransistorNmos: 1.42551e+07 muA
** DiodeTransistorPmos: -1.72606e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.23301  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 4.25  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.784001  V
** outVoltageBiasXXnXX0: 0.769001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40001  V
** innerTransistorStack1Load1: 0.228001  V
** innerTransistorStack2Load1: 0.228001  V
** sourceTransconductance: 3.21801  V
** innerStageBias: 4.48901  V
** innerTransconductance: 0.212001  V
** inner: 4.40001  V
** inner: 0.212001  V


.END