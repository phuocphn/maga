** Name: two_stage_single_output_op_amp_53_8

.MACRO two_stage_single_output_op_amp_53_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=8e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=132e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=10e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=488e-6
mSecondStage1StageBias12 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=475e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=8e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=87e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=555e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=87e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=115e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=218e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_53_8

** Expected Performance Values: 
** Gain: 118 dB
** Power consumption: 6.31901 mW
** Area: 8239 (mu_m)^2
** Transit frequency: 3.24101 MHz
** Transit frequency with error factor: 3.24074 MHz
** Slew rate: 7.7623 V/mu_s
** Phase margin: 69.328°
** CMRR: 133 dB
** VoutMax: 4.25 V
** VoutMin: 0.480001 V
** VcmMax: 5.17001 V
** VcmMin: 1.07001 V


** Expected Currents: 
** NormalTransistorPmos: -1.16595e+08 muA
** NormalTransistorPmos: -2.16839e+08 muA
** NormalTransistorPmos: -3.51479e+07 muA
** NormalTransistorPmos: -5.27209e+07 muA
** NormalTransistorPmos: -3.51479e+07 muA
** NormalTransistorPmos: -5.27209e+07 muA
** DiodeTransistorNmos: 3.51471e+07 muA
** DiodeTransistorNmos: 3.51461e+07 muA
** NormalTransistorNmos: 3.51471e+07 muA
** NormalTransistorNmos: 3.51461e+07 muA
** NormalTransistorNmos: 3.51471e+07 muA
** NormalTransistorNmos: 1.75741e+07 muA
** NormalTransistorNmos: 1.75741e+07 muA
** NormalTransistorNmos: 8.0502e+08 muA
** NormalTransistorNmos: 8.05019e+08 muA
** NormalTransistorPmos: -8.05019e+08 muA
** DiodeTransistorNmos: 1.16596e+08 muA
** DiodeTransistorNmos: 2.1684e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.08501  V
** outVoltageBiasXXnXX2: 0.685001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.776001  V
** innerTransistorStack2Load2: 0.774001  V
** out1: 1.50201  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.71201  V
** innerStageBias: 0.480001  V


.END