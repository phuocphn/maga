** Name: two_stage_single_output_op_amp_160_1

.MACRO two_stage_single_output_op_amp_160_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=28e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=7e-6
mMainBias3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=203e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mSimpleFirstStageLoad6 FirstStageYout1 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=40e-6
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad8 outFirstStage ibias sourceNmos sourceNmos nmos4 L=6e-6 W=40e-6
mMainBias9 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=302e-6
mMainBias10 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=430e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=101e-6
mSimpleFirstStageLoad12 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=7e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=43e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=203e-6
mSecondStage1StageBias15 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=227e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=9e-6 W=9e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=101e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.30001e-12
.EOM two_stage_single_output_op_amp_160_1

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 12.9851 mW
** Area: 7563 (mu_m)^2
** Transit frequency: 3.20001 MHz
** Transit frequency with error factor: 3.19999 MHz
** Slew rate: 3.54838 V/mu_s
** Phase margin: 60.1606°
** CMRR: 79 dB
** VoutMax: 4.25 V
** VoutMin: 0.210001 V
** VcmMax: 3.35001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorNmos: 1.0665e+08 muA
** NormalTransistorNmos: 1.52301e+08 muA
** NormalTransistorPmos: -2.88799e+06 muA
** NormalTransistorPmos: -2.88799e+06 muA
** DiodeTransistorPmos: -2.88799e+06 muA
** NormalTransistorNmos: 1.41261e+07 muA
** NormalTransistorNmos: 1.41261e+07 muA
** NormalTransistorPmos: -2.24789e+07 muA
** DiodeTransistorPmos: -2.24799e+07 muA
** NormalTransistorPmos: -1.12389e+07 muA
** NormalTransistorPmos: -1.12389e+07 muA
** NormalTransistorNmos: 2.29977e+09 muA
** NormalTransistorPmos: -2.29976e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.06649e+08 muA
** NormalTransistorPmos: -1.0665e+08 muA
** DiodeTransistorPmos: -1.523e+08 muA


** Expected Voltages: 
** ibias: 0.564001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.617001  V
** outInputVoltageBiasXXpXX1: 3.53001  V
** outSourceVoltageBiasXXpXX1: 4.26501  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.03201  V
** out1: 3.06401  V
** sourceTransconductance: 3.24001  V
** inner: 4.26501  V


.END