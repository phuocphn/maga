** Name: two_stage_single_output_op_amp_79_6

.MACRO two_stage_single_output_op_amp_79_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=15e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=19e-6
mMainBias3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=21e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=14e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=525e-6
mMainBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=197e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=101e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=101e-6
mFoldedCascodeFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=345e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=345e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=68e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=110e-6
mMainBias15 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=321e-6
mSecondStage1Transconductor16 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=574e-6
mFoldedCascodeFirstStageLoad17 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=39e-6
mMainBias18 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=44e-6
mFoldedCascodeFirstStageLoad19 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=239e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mMainBias22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=14e-6
mSecondStage1StageBias23 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=525e-6
mFoldedCascodeFirstStageLoad24 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=239e-6
mMainBias25 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=48e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.6001e-12
.EOM two_stage_single_output_op_amp_79_6

** Expected Performance Values: 
** Gain: 176 dB
** Power consumption: 10.7891 mW
** Area: 14872 (mu_m)^2
** Transit frequency: 6.74801 MHz
** Transit frequency with error factor: 6.74827 MHz
** Slew rate: 4.68203 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 3.25 V
** VoutMin: 0.490001 V
** VcmMax: 4.66001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 2.91311e+07 muA
** NormalTransistorNmos: 2.13221e+08 muA
** NormalTransistorPmos: -4.87362e+08 muA
** NormalTransistorPmos: -9.67449e+07 muA
** NormalTransistorPmos: -1.62453e+08 muA
** NormalTransistorPmos: -9.67449e+07 muA
** NormalTransistorPmos: -1.62453e+08 muA
** NormalTransistorNmos: 9.67441e+07 muA
** NormalTransistorNmos: 9.67431e+07 muA
** NormalTransistorNmos: 9.67441e+07 muA
** NormalTransistorNmos: 9.67431e+07 muA
** NormalTransistorNmos: 1.3142e+08 muA
** NormalTransistorNmos: 1.31419e+08 muA
** NormalTransistorNmos: 6.57101e+07 muA
** NormalTransistorNmos: 6.57101e+07 muA
** NormalTransistorNmos: 1.09326e+09 muA
** NormalTransistorNmos: 1.09326e+09 muA
** NormalTransistorPmos: -1.09325e+09 muA
** DiodeTransistorPmos: -1.09325e+09 muA
** DiodeTransistorNmos: 4.87363e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.91319e+07 muA
** NormalTransistorPmos: -2.91329e+07 muA
** DiodeTransistorPmos: -2.1322e+08 muA
** DiodeTransistorPmos: -2.1322e+08 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.749001  V
** outInputVoltageBiasXXpXX1: 2.68401  V
** outSourceVoltageBiasXXpXX1: 3.84201  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX1: 0.954001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.398001  V
** innerTransistorStack1Load2: 0.377001  V
** innerTransistorStack2Load2: 0.377001  V
** out1: 0.555001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 0.399001  V
** inner: 3.83701  V


.END