** Name: two_stage_single_output_op_amp_75_6

.MACRO two_stage_single_output_op_amp_75_6 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=126e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=5e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=491e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=234e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=126e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=227e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=227e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=94e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mMainBias14 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=82e-6
mSecondStage1Transconductor15 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=596e-6
mFoldedCascodeFirstStageLoad16 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=63e-6
mMainBias17 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=15e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=591e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=38e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=38e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=491e-6
mFoldedCascodeFirstStageLoad23 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=591e-6
mMainBias24 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.3001e-12
.EOM two_stage_single_output_op_amp_75_6

** Expected Performance Values: 
** Gain: 179 dB
** Power consumption: 14.9911 mW
** Area: 6944 (mu_m)^2
** Transit frequency: 15.7301 MHz
** Transit frequency with error factor: 15.7302 MHz
** Slew rate: 12.3459 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 3.14001 V
** VoutMin: 0.380001 V
** VcmMax: 4.66001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorNmos: 1.86291e+07 muA
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -2.70062e+08 muA
** NormalTransistorPmos: -2.40025e+08 muA
** NormalTransistorPmos: -3.84143e+08 muA
** NormalTransistorPmos: -2.40025e+08 muA
** NormalTransistorPmos: -3.84143e+08 muA
** DiodeTransistorNmos: 2.40026e+08 muA
** NormalTransistorNmos: 2.40026e+08 muA
** NormalTransistorNmos: 2.40026e+08 muA
** NormalTransistorNmos: 2.88234e+08 muA
** NormalTransistorNmos: 2.88233e+08 muA
** NormalTransistorNmos: 1.44118e+08 muA
** NormalTransistorNmos: 1.44118e+08 muA
** NormalTransistorNmos: 1.82968e+09 muA
** NormalTransistorNmos: 1.82968e+09 muA
** NormalTransistorPmos: -1.82967e+09 muA
** DiodeTransistorPmos: -1.82967e+09 muA
** DiodeTransistorNmos: 2.70063e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.86299e+07 muA
** NormalTransistorPmos: -1.86309e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.594001  V
** outInputVoltageBiasXXpXX1: 2.57401  V
** outSourceVoltageBiasXXpXX1: 3.78701  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX1: 0.967001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.371001  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 0.371001  V
** inner: 3.78101  V


.END