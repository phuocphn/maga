** Name: two_stage_single_output_op_amp_13_7

.MACRO two_stage_single_output_op_amp_13_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=36e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=5e-6 W=36e-6
mSimpleFirstStageTransconductor4 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=11e-6
mSimpleFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mSecondStage1StageBias6 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=271e-6
mSimpleFirstStageTransconductor7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=11e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=36e-6
mSecondStage1Transconductor9 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=36e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_13_7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 2.43201 mW
** Area: 1696 (mu_m)^2
** Transit frequency: 2.75801 MHz
** Transit frequency with error factor: 2.75362 MHz
** Slew rate: 6.55136 V/mu_s
** Phase margin: 61.3065°
** CMRR: 95 dB
** negPSRR: 93 dB
** posPSRR: 86 dB
** VoutMax: 4.25 V
** VoutMin: 0.200001 V
** VcmMax: 3.54001 V
** VcmMin: 0.980001 V


** Expected Currents: 
** DiodeTransistorPmos: -1.47869e+07 muA
** NormalTransistorPmos: -1.47879e+07 muA
** NormalTransistorPmos: -1.47869e+07 muA
** DiodeTransistorPmos: -1.47879e+07 muA
** NormalTransistorNmos: 2.95721e+07 muA
** NormalTransistorNmos: 1.47861e+07 muA
** NormalTransistorNmos: 1.47861e+07 muA
** NormalTransistorNmos: 4.46749e+08 muA
** NormalTransistorPmos: -4.46748e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.03401  V
** innerTransistorStack1Load1: 4.03401  V
** out1: 3.13201  V
** sourceTransconductance: 1.71601  V


.END