** Name: two_stage_single_output_op_amp_137_6

.MACRO two_stage_single_output_op_amp_137_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=55e-6
mSecondStage1StageBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=23e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=5e-6 W=29e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=29e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=22e-6
mMainBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=109e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=358e-6
mSimpleFirstStageLoad8 FirstStageYinnerOutputLoad1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=29e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=163e-6
mMainBias10 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mSecondStage1Transconductor11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=245e-6
mSimpleFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=29e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=33e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=29e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=122e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=109e-6
mMainBias17 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=357e-6
mSecondStage1StageBias18 out inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=358e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=29e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=33e-6
mMainBias21 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=111e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_137_6

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 3.05401 mW
** Area: 11141 (mu_m)^2
** Transit frequency: 2.86901 MHz
** Transit frequency with error factor: 2.84692 MHz
** Slew rate: 6.30073 V/mu_s
** Phase margin: 61.3065°
** CMRR: 75 dB
** VoutMax: 3.61001 V
** VoutMin: 0.320001 V
** VcmMax: 3.47001 V
** VcmMin: -0.379999 V


** Expected Currents: 
** NormalTransistorNmos: 4.73961e+07 muA
** NormalTransistorPmos: -5.12439e+07 muA
** NormalTransistorPmos: -1.62924e+08 muA
** DiodeTransistorPmos: -5.88889e+07 muA
** NormalTransistorPmos: -5.88889e+07 muA
** NormalTransistorPmos: -5.88889e+07 muA
** DiodeTransistorPmos: -5.88889e+07 muA
** NormalTransistorNmos: 8.70501e+07 muA
** NormalTransistorNmos: 8.70501e+07 muA
** NormalTransistorPmos: -5.63229e+07 muA
** NormalTransistorPmos: -2.81619e+07 muA
** NormalTransistorPmos: -2.81619e+07 muA
** NormalTransistorNmos: 1.55227e+08 muA
** NormalTransistorNmos: 1.55228e+08 muA
** NormalTransistorPmos: -1.55226e+08 muA
** DiodeTransistorPmos: -1.55227e+08 muA
** DiodeTransistorNmos: 5.12431e+07 muA
** DiodeTransistorNmos: 1.62925e+08 muA
** DiodeTransistorPmos: -4.73969e+07 muA
** NormalTransistorPmos: -4.73979e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.15901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.593001  V
** inputVoltageBiasXXpXX1: 3.04401  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.02201  V
** outVoltageBiasXXnXX1: 0.728001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerSourceLoad1: 3.68601  V
** innerTransistorStack1Load1: 3.68601  V
** sourceTransconductance: 3.75201  V
** innerTransconductance: 0.150001  V
** inner: 4.01901  V


.END