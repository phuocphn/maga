** Name: two_stage_single_output_op_amp_64_1

.MACRO two_stage_single_output_op_amp_64_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=21e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=9e-6 W=129e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=9e-6 W=118e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=11e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=74e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=29e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=71e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=71e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=57e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=29e-6
mMainBias13 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mMainBias14 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=47e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=9e-6 W=129e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=74e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=11e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=536e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=9e-6 W=118e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_64_1

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 3.61701 mW
** Area: 6988 (mu_m)^2
** Transit frequency: 3.58801 MHz
** Transit frequency with error factor: 3.5877 MHz
** Slew rate: 3.95386 V/mu_s
** Phase margin: 67.0361°
** CMRR: 139 dB
** VoutMax: 4.74001 V
** VoutMin: 0.520001 V
** VcmMax: 3.36001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.68001e+06 muA
** NormalTransistorNmos: 1.80841e+07 muA
** NormalTransistorNmos: 1.79201e+07 muA
** NormalTransistorNmos: 2.70461e+07 muA
** NormalTransistorNmos: 1.79201e+07 muA
** NormalTransistorNmos: 2.70461e+07 muA
** DiodeTransistorPmos: -1.79209e+07 muA
** DiodeTransistorPmos: -1.79219e+07 muA
** NormalTransistorPmos: -1.79209e+07 muA
** NormalTransistorPmos: -1.79219e+07 muA
** NormalTransistorPmos: -1.82549e+07 muA
** DiodeTransistorPmos: -1.82559e+07 muA
** NormalTransistorPmos: -9.12699e+06 muA
** NormalTransistorPmos: -9.12699e+06 muA
** NormalTransistorNmos: 6.38458e+08 muA
** NormalTransistorPmos: -6.38457e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.68099e+06 muA
** NormalTransistorPmos: -2.68199e+06 muA
** DiodeTransistorPmos: -1.80849e+07 muA


** Expected Voltages: 
** ibias: 1.12701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.922001  V
** outInputVoltageBiasXXpXX1: 3.54001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.27001  V
** outVoltageBiasXXpXX2: 4.17701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.17101  V
** innerTransistorStack2Load2: 4.17001  V
** out1: 3.33001  V
** sourceGCC1: 0.530001  V
** sourceGCC2: 0.530001  V
** sourceTransconductance: 3.24201  V
** inner: 4.26901  V


.END