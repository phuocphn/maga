** Name: two_stage_single_output_op_amp_68_1

.MACRO two_stage_single_output_op_amp_68_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=5e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=39e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=16e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=73e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=7e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=256e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=7e-6
mMainBias13 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias14 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=103e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=103e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=73e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=16e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=596e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=39e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_68_1

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 6.23501 mW
** Area: 6527 (mu_m)^2
** Transit frequency: 3.66601 MHz
** Transit frequency with error factor: 3.66624 MHz
** Slew rate: 3.85123 V/mu_s
** Phase margin: 76.2034°
** CMRR: 142 dB
** VoutMax: 4.33001 V
** VoutMin: 0.620001 V
** VcmMax: 3.30001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.92401e+06 muA
** NormalTransistorNmos: 1.00071e+07 muA
** NormalTransistorNmos: 1.73671e+07 muA
** NormalTransistorNmos: 2.61601e+07 muA
** NormalTransistorNmos: 1.73671e+07 muA
** NormalTransistorNmos: 2.61601e+07 muA
** DiodeTransistorPmos: -1.73679e+07 muA
** NormalTransistorPmos: -1.73689e+07 muA
** NormalTransistorPmos: -1.73679e+07 muA
** DiodeTransistorPmos: -1.73689e+07 muA
** NormalTransistorPmos: -1.75889e+07 muA
** DiodeTransistorPmos: -1.75899e+07 muA
** NormalTransistorPmos: -8.79399e+06 muA
** NormalTransistorPmos: -8.79399e+06 muA
** NormalTransistorNmos: 1.17065e+09 muA
** NormalTransistorPmos: -1.17064e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.92499e+06 muA
** NormalTransistorPmos: -3.92599e+06 muA
** DiodeTransistorPmos: -1.00079e+07 muA


** Expected Voltages: 
** ibias: 1.22801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 1.02301  V
** outInputVoltageBiasXXpXX1: 3.46801  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.23401  V
** outVoltageBiasXXpXX2: 3.77001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.27801  V
** innerTransistorStack2Load2: 4.27801  V
** out1: 3.55601  V
** sourceGCC1: 0.525001  V
** sourceGCC2: 0.525001  V
** sourceTransconductance: 3.23301  V
** inner: 4.23401  V


.END