** Name: one_stage_single_output_op_amp116

.MACRO one_stage_single_output_op_amp116 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=13e-6
mTelescopicFirstStageStageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=133e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=27e-6
mTelescopicFirstStageLoad4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=29e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
mTelescopicFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=52e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=13e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=13e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mMainBias10 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mTelescopicFirstStageLoad11 out outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=52e-6
mTelescopicFirstStageStageBias12 sourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=133e-6
mTelescopicFirstStageLoad13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=29e-6
mTelescopicFirstStageLoad14 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=26e-6
mMainBias15 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=40e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp116

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 0.595001 mW
** Area: 1874 (mu_m)^2
** Transit frequency: 2.62401 MHz
** Transit frequency with error factor: 2.62371 MHz
** Slew rate: 5.05122 V/mu_s
** Phase margin: 87.6626°
** CMRR: 145 dB
** VoutMax: 3.89001 V
** VoutMin: 1.03001 V
** VcmMax: 4.15001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 7.75901e+06 muA
** NormalTransistorPmos: -5.16359e+07 muA
** NormalTransistorNmos: 2.47621e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorPmos: -2.47629e+07 muA
** NormalTransistorPmos: -2.47619e+07 muA
** DiodeTransistorPmos: -2.47629e+07 muA
** NormalTransistorNmos: 1.01159e+08 muA
** DiodeTransistorNmos: 1.0116e+08 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 5.16351e+07 muA
** DiodeTransistorPmos: -7.75999e+06 muA


** Expected Voltages: 
** ibias: 1.13901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.77501  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.570001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.12601  V
** out1: 3.33001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.569001  V


.END