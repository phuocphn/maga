** Name: symmetrical_op_amp118

.MACRO symmetrical_op_amp118 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=11e-6
mSecondStage1StageBias2 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=47e-6
mSymmetricalFirstStageTransconductor5 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=33e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias7 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos4 L=1e-6 W=25e-6
mSymmetricalFirstStageTransconductor8 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=33e-6
mMainBias9 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=7e-6 W=111e-6
mSymmetricalFirstStageLoad10 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=13e-6
mSymmetricalFirstStageLoad11 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=13e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=31e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor13 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=31e-6
mSymmetricalFirstStageLoad14 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=52e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=125e-6
mSecondStage1Transconductor16 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=125e-6
mSymmetricalFirstStageLoad17 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=52e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp118

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 1.26901 mW
** Area: 2558 (mu_m)^2
** Transit frequency: 3.05701 MHz
** Transit frequency with error factor: 3.05686 MHz
** Slew rate: 5.02775 V/mu_s
** Phase margin: 85.9437°
** CMRR: 140 dB
** negPSRR: 128 dB
** posPSRR: 61 dB
** VoutMax: 4.25 V
** VoutMin: 0.900001 V
** VcmMax: 4.81001 V
** VcmMin: 0.940001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01052e+08 muA
** NormalTransistorPmos: -2.09709e+07 muA
** NormalTransistorPmos: -2.09719e+07 muA
** NormalTransistorPmos: -2.09709e+07 muA
** NormalTransistorPmos: -2.09719e+07 muA
** NormalTransistorNmos: 4.19411e+07 muA
** NormalTransistorNmos: 2.09701e+07 muA
** NormalTransistorNmos: 2.09701e+07 muA
** NormalTransistorNmos: 5.03601e+07 muA
** DiodeTransistorNmos: 5.03591e+07 muA
** NormalTransistorPmos: -5.03609e+07 muA
** NormalTransistorPmos: -5.03599e+07 muA
** NormalTransistorNmos: 5.03601e+07 muA
** NormalTransistorPmos: -5.03609e+07 muA
** NormalTransistorPmos: -5.03599e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.01051e+08 muA


** Expected Voltages: 
** ibias: 0.678001  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** inStageBiasComplementarySecondStage: 0.749001  V
** innerComplementarySecondStage: 1.30801  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.83401  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END