** Name: two_stage_single_output_op_amp_33_11

.MACRO two_stage_single_output_op_amp_33_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=9e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=275e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=109e-6
mSimpleFirstStageTransconductor5 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=21e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=29e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=391e-6
mSecondStage1StageBias9 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=250e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=21e-6
mMainBias11 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=139e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=275e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=480e-6
mSecondStage1Transconductor14 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=8e-6 W=600e-6
mSimpleFirstStageLoad15 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=8e-6 W=271e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.20001e-12
.EOM two_stage_single_output_op_amp_33_11

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 2.84101 mW
** Area: 14646 (mu_m)^2
** Transit frequency: 2.77501 MHz
** Transit frequency with error factor: 2.77456 MHz
** Slew rate: 3.54781 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** negPSRR: 99 dB
** posPSRR: 94 dB
** VoutMax: 4.25 V
** VoutMin: 0.75 V
** VcmMax: 4.53001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorNmos: 1.3834e+08 muA
** DiodeTransistorPmos: -1.47149e+07 muA
** NormalTransistorPmos: -1.47149e+07 muA
** NormalTransistorPmos: -1.47149e+07 muA
** NormalTransistorNmos: 2.94291e+07 muA
** NormalTransistorNmos: 2.94301e+07 muA
** NormalTransistorNmos: 1.47141e+07 muA
** NormalTransistorNmos: 1.47141e+07 muA
** NormalTransistorNmos: 3.9039e+08 muA
** NormalTransistorNmos: 3.90389e+08 muA
** NormalTransistorPmos: -3.90389e+08 muA
** NormalTransistorPmos: -3.9039e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.38339e+08 muA


** Expected Voltages: 
** ibias: 1.125  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.22301  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.28101  V
** innerStageBias: 0.565001  V
** innerTransistorStack2Load1: 4.40601  V
** sourceTransconductance: 1.89101  V
** innerStageBias: 0.527001  V
** innerTransconductance: 4.78701  V


.END