** Name: one_stage_single_output_op_amp101

.MACRO one_stage_single_output_op_amp101 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=21e-6
mMainBias4 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=8e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mTelescopicFirstStageLoad7 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=30e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=42e-6
mTelescopicFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=234e-6
mTelescopicFirstStageLoad10 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=65e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=130e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=130e-6
mTelescopicFirstStageLoad13 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=65e-6
mMainBias14 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=589e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp101

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 1.34101 mW
** Area: 3097 (mu_m)^2
** Transit frequency: 3 MHz
** Transit frequency with error factor: 2.99972 MHz
** Slew rate: 11.8321 V/mu_s
** Phase margin: 87.6626°
** CMRR: 133 dB
** VoutMax: 3.08001 V
** VoutMin: 0.890001 V
** VcmMax: 3 V
** VcmMin: 0.820001 V


** Expected Currents: 
** NormalTransistorNmos: 5.29661e+07 muA
** NormalTransistorPmos: -1.11519e+07 muA
** NormalTransistorPmos: -9.19949e+07 muA
** NormalTransistorPmos: -9.19959e+07 muA
** NormalTransistorNmos: 9.19941e+07 muA
** NormalTransistorNmos: 9.19951e+07 muA
** DiodeTransistorNmos: 9.19941e+07 muA
** NormalTransistorPmos: -2.36957e+08 muA
** NormalTransistorPmos: -2.36958e+08 muA
** NormalTransistorPmos: -9.19949e+07 muA
** NormalTransistorPmos: -9.19949e+07 muA
** DiodeTransistorNmos: 1.11511e+07 muA
** DiodeTransistorPmos: -5.29669e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.648001  V
** outVoltageBiasXXpXX1: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.54901  V
** innerSourceLoad2: 0.705001  V
** innerStageBias: 4.18501  V
** out1: 1.30001  V
** sourceGCC1: 2.98801  V
** sourceGCC2: 2.98801  V


.END