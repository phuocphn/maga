** Name: one_stage_single_output_op_amp105

.MACRO one_stage_single_output_op_amp105 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=16e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=30e-6
mMainBias5 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=16e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
mTelescopicFirstStageLoad8 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=16e-6
mMainBias9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mTelescopicFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=56e-6
mTelescopicFirstStageLoad11 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=68e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=237e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=237e-6
mTelescopicFirstStageLoad14 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=68e-6
mMainBias15 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=11e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=562e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp105

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 0.782001 mW
** Area: 5326 (mu_m)^2
** Transit frequency: 2.78501 MHz
** Transit frequency with error factor: 2.78549 MHz
** Slew rate: 5.69493 V/mu_s
** Phase margin: 78.4953°
** CMRR: 139 dB
** VoutMax: 3.07001 V
** VoutMin: 0.75 V
** VcmMax: 3 V
** VcmMin: 1.09001 V


** Expected Currents: 
** NormalTransistorNmos: 2.70371e+07 muA
** NormalTransistorPmos: -2.23989e+07 muA
** NormalTransistorPmos: -4.35e+07 muA
** NormalTransistorPmos: -4.35e+07 muA
** DiodeTransistorNmos: 4.34991e+07 muA
** DiodeTransistorNmos: 4.34981e+07 muA
** NormalTransistorNmos: 4.34991e+07 muA
** NormalTransistorNmos: 4.34981e+07 muA
** NormalTransistorPmos: -1.14034e+08 muA
** NormalTransistorPmos: -1.14033e+08 muA
** NormalTransistorPmos: -4.34989e+07 muA
** NormalTransistorPmos: -4.34989e+07 muA
** DiodeTransistorNmos: 2.23981e+07 muA
** DiodeTransistorPmos: -2.70379e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.20301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX2: 3.96101  V
** outVoltageBiasXXnXX0: 0.568001  V
** outVoltageBiasXXpXX1: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.31101  V
** innerStageBias: 3.91701  V
** innerTransistorStack1Load2: 0.574001  V
** innerTransistorStack2Load2: 0.573001  V
** out1: 1.15801  V
** sourceGCC1: 2.99901  V
** sourceGCC2: 2.99901  V


.END