** Name: symmetrical_op_amp35

.MACRO symmetrical_op_amp35 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=11e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=11e-6
mSymmetricalFirstStageLoad4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=90e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=119e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=24e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=24e-6
mMainBias12 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=94e-6
mSymmetricalFirstStageStageBias13 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=207e-6
mSymmetricalFirstStageStageBias14 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=83e-6
mSecondStage1StageBias15 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=119e-6
mMainBias16 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=6e-6 W=507e-6
mSymmetricalFirstStageTransconductor17 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=107e-6
mMainBias18 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=27e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=12e-6
mSymmetricalFirstStageTransconductor20 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=107e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp35

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 0.988001 mW
** Area: 8042 (mu_m)^2
** Transit frequency: 3.54001 MHz
** Transit frequency with error factor: 3.53978 MHz
** Slew rate: 3.50003 V/mu_s
** Phase margin: 81.933°
** CMRR: 139 dB
** negPSRR: 54 dB
** posPSRR: 71 dB
** VoutMax: 4.25 V
** VoutMin: 0.610001 V
** VcmMax: 3.35001 V
** VcmMin: 0.130001 V


** Expected Currents: 
** NormalTransistorNmos: 2.53821e+07 muA
** NormalTransistorPmos: -3.01399e+06 muA
** NormalTransistorPmos: -5.66159e+07 muA
** DiodeTransistorNmos: 1.15061e+07 muA
** DiodeTransistorNmos: 1.15061e+07 muA
** NormalTransistorPmos: -2.30149e+07 muA
** NormalTransistorPmos: -2.30159e+07 muA
** NormalTransistorPmos: -1.15069e+07 muA
** NormalTransistorPmos: -1.15069e+07 muA
** NormalTransistorNmos: 3.50131e+07 muA
** NormalTransistorNmos: 3.50121e+07 muA
** NormalTransistorPmos: -3.50139e+07 muA
** NormalTransistorPmos: -3.50149e+07 muA
** DiodeTransistorPmos: -3.45179e+07 muA
** NormalTransistorNmos: 3.45171e+07 muA
** NormalTransistorNmos: 3.45181e+07 muA
** DiodeTransistorNmos: 3.01301e+06 muA
** DiodeTransistorNmos: 5.66151e+07 muA
** DiodeTransistorPmos: -2.53829e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 1.01201  V
** inSourceTransconductanceComplementarySecondStage: 0.692001  V
** innerComplementarySecondStage: 4.25501  V
** inputVoltageBiasXXnXX0: 0.584001  V
** out: 2.5  V
** outFirstStage: 0.692001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.42601  V
** sourceTransconductance: 3.21901  V
** innerStageBias: 4.81901  V
** innerTransconductance: 0.287001  V
** inner: 0.287001  V


.END