** Name: two_stage_single_output_op_amp_190_12

.MACRO two_stage_single_output_op_amp_190_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=7e-6 W=37e-6
mMainBias2 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=8e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=161e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=34e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=372e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=126e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=299e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=33e-6
mSimpleFirstStageLoad9 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=7e-6 W=37e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=34e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=161e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mSecondStage1StageBias13 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=372e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=30e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=33e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=256e-6
mMainBias17 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=98e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=517e-6
mSimpleFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=517e-6
mSimpleFirstStageLoad20 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=128e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=531e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=503e-6
mSimpleFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=128e-6
mMainBias24 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=290e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5e-12
.EOM two_stage_single_output_op_amp_190_12

** Expected Performance Values: 
** Gain: 144 dB
** Power consumption: 7.17301 mW
** Area: 13098 (mu_m)^2
** Transit frequency: 5.28301 MHz
** Transit frequency with error factor: 5.28026 MHz
** Slew rate: 4.97875 V/mu_s
** Phase margin: 60.1606°
** CMRR: 119 dB
** VoutMax: 4.33001 V
** VoutMin: 0.890001 V
** VcmMax: 4.66001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 3.14136e+08 muA
** NormalTransistorNmos: 1.20256e+08 muA
** NormalTransistorPmos: -1.17778e+08 muA
** NormalTransistorNmos: 1.9537e+08 muA
** NormalTransistorNmos: 1.9537e+08 muA
** DiodeTransistorNmos: 1.9537e+08 muA
** NormalTransistorPmos: -2.0794e+08 muA
** NormalTransistorPmos: -2.07941e+08 muA
** NormalTransistorPmos: -2.0794e+08 muA
** NormalTransistorPmos: -2.07941e+08 muA
** NormalTransistorNmos: 2.51411e+07 muA
** DiodeTransistorNmos: 2.51401e+07 muA
** NormalTransistorNmos: 1.25711e+07 muA
** NormalTransistorNmos: 1.25711e+07 muA
** NormalTransistorNmos: 4.56478e+08 muA
** DiodeTransistorNmos: 4.56479e+08 muA
** NormalTransistorPmos: -4.56477e+08 muA
** NormalTransistorPmos: -4.56478e+08 muA
** DiodeTransistorNmos: 1.17779e+08 muA
** NormalTransistorNmos: 1.17778e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.14135e+08 muA
** DiodeTransistorPmos: -1.20255e+08 muA


** Expected Voltages: 
** ibias: 1.29201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.21601  V
** outInputVoltageBiasXXnXX1: 1.22601  V
** outSourceVoltageBiasXXnXX1: 0.613001  V
** outSourceVoltageBiasXXnXX2: 0.647001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.28601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.85001  V
** innerTransistorStack2Load1: 1.06701  V
** innerTransistorStack2Load2: 4.85001  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.69901  V
** inner: 0.613001  V
** inner: 0.643001  V


.END