** Name: two_stage_single_output_op_amp_24_4

.MACRO two_stage_single_output_op_amp_24_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=59e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=8e-6 W=51e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=88e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=122e-6
mMainBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
mSimpleFirstStageLoad7 FirstStageYinnerSourceLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=53e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=92e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=92e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=268e-6
mSecondStage1Transconductor11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=357e-6
mSimpleFirstStageLoad12 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=53e-6
mMainBias13 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=194e-6
mSimpleFirstStageTransconductor14 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=57e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=122e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=135e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=88e-6
mSecondStage1StageBias18 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=8e-6 W=600e-6
mSimpleFirstStageTransconductor19 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=57e-6
mMainBias20 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=9e-6
mMainBias21 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=18e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.3001e-12
.EOM two_stage_single_output_op_amp_24_4

** Expected Performance Values: 
** Gain: 147 dB
** Power consumption: 1.56201 mW
** Area: 14998 (mu_m)^2
** Transit frequency: 2.92901 MHz
** Transit frequency with error factor: 2.92661 MHz
** Slew rate: 4.10073 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** negPSRR: 105 dB
** posPSRR: 172 dB
** VoutMax: 3.33001 V
** VoutMin: 0.300001 V
** VcmMax: 3.04001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.70741e+07 muA
** NormalTransistorPmos: -1.14219e+07 muA
** NormalTransistorPmos: -2.28449e+07 muA
** NormalTransistorNmos: 2.52831e+07 muA
** NormalTransistorNmos: 2.52821e+07 muA
** NormalTransistorNmos: 2.52831e+07 muA
** NormalTransistorNmos: 2.52821e+07 muA
** NormalTransistorPmos: -5.05689e+07 muA
** DiodeTransistorPmos: -5.05699e+07 muA
** NormalTransistorPmos: -2.52839e+07 muA
** NormalTransistorPmos: -2.52839e+07 muA
** NormalTransistorNmos: 1.70447e+08 muA
** NormalTransistorNmos: 1.70446e+08 muA
** NormalTransistorPmos: -1.70446e+08 muA
** NormalTransistorPmos: -1.70447e+08 muA
** DiodeTransistorNmos: 1.14211e+07 muA
** DiodeTransistorNmos: 2.28441e+07 muA
** DiodeTransistorPmos: -3.70749e+07 muA
** NormalTransistorPmos: -3.70759e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.82501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.26001  V
** outSourceVoltageBiasXXpXX1: 4.13001  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX0: 0.556001  V
** outVoltageBiasXXnXX1: 0.705001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.28601  V
** innerStageBias: 3.74401  V
** innerTransconductance: 0.150001  V
** inner: 4.13001  V


.END