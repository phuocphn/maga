** Name: two_stage_single_output_op_amp_12_8

.MACRO two_stage_single_output_op_amp_12_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=30e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
mMainBias3 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=15e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSimpleFirstStageTransconductor5 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=18e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=6e-6 W=105e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=600e-6
mSecondStage1StageBias8 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=6e-6 W=83e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=18e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=30e-6
mMainBias11 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=30e-6
mSimpleFirstStageLoad12 FirstStageYinnerSourceLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=4e-6 W=150e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=48e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=48e-6
mMainBias15 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=139e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=368e-6
mSimpleFirstStageLoad17 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=150e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9e-12
.EOM two_stage_single_output_op_amp_12_8

** Expected Performance Values: 
** Gain: 107 dB
** Power consumption: 1.77501 mW
** Area: 8872 (mu_m)^2
** Transit frequency: 4.02001 MHz
** Transit frequency with error factor: 4.01806 MHz
** Slew rate: 3.79203 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** negPSRR: 130 dB
** posPSRR: 107 dB
** VoutMax: 4.83001 V
** VoutMin: 0.560001 V
** VcmMax: 5.16001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorNmos: 9.97501e+06 muA
** NormalTransistorNmos: 9.85601e+06 muA
** NormalTransistorPmos: -9.07599e+07 muA
** NormalTransistorPmos: -1.71679e+07 muA
** NormalTransistorPmos: -1.71689e+07 muA
** NormalTransistorPmos: -1.71679e+07 muA
** NormalTransistorPmos: -1.71689e+07 muA
** NormalTransistorNmos: 3.43351e+07 muA
** NormalTransistorNmos: 1.71671e+07 muA
** NormalTransistorNmos: 1.71671e+07 muA
** NormalTransistorNmos: 2.0016e+08 muA
** NormalTransistorNmos: 2.00159e+08 muA
** NormalTransistorPmos: -2.00159e+08 muA
** DiodeTransistorNmos: 9.07591e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.97599e+06 muA
** DiodeTransistorPmos: -9.85699e+06 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.970001  V
** out: 2.5  V
** outFirstStage: 4.26101  V
** outVoltageBiasXXpXX0: 3.82901  V
** outVoltageBiasXXpXX1: 3.69701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.19001  V
** innerTransistorStack1Load1: 4.42101  V
** innerTransistorStack2Load1: 4.42101  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.153001  V


.END