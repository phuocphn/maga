** Name: two_stage_single_output_op_amp_77_11

.MACRO two_stage_single_output_op_amp_77_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=24e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=5e-6 W=24e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=13e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=302e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=78e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=27e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=5e-6 W=24e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=8e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=8e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=13e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=534e-6
mMainBias13 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=60e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=559e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=24e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=299e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerOutputLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=57e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=203e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=203e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=570e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=278e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=57e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_77_11

** Expected Performance Values: 
** Gain: 172 dB
** Power consumption: 3.27601 mW
** Area: 11094 (mu_m)^2
** Transit frequency: 2.72101 MHz
** Transit frequency with error factor: 2.72081 MHz
** Slew rate: 3.90398 V/mu_s
** Phase margin: 67.6091°
** CMRR: 138 dB
** VoutMax: 4.28001 V
** VoutMin: 0.710001 V
** VcmMax: 5.21001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorNmos: 1.97991e+08 muA
** NormalTransistorNmos: 3.93381e+07 muA
** NormalTransistorPmos: -1.76569e+07 muA
** NormalTransistorPmos: -2.64839e+07 muA
** NormalTransistorPmos: -1.76609e+07 muA
** NormalTransistorPmos: -2.64899e+07 muA
** DiodeTransistorNmos: 1.76581e+07 muA
** DiodeTransistorNmos: 1.76591e+07 muA
** NormalTransistorNmos: 1.76601e+07 muA
** NormalTransistorNmos: 1.76591e+07 muA
** NormalTransistorNmos: 1.76571e+07 muA
** NormalTransistorNmos: 1.76581e+07 muA
** NormalTransistorNmos: 8.82801e+06 muA
** NormalTransistorNmos: 8.82801e+06 muA
** NormalTransistorNmos: 3.54897e+08 muA
** NormalTransistorNmos: 3.54896e+08 muA
** NormalTransistorPmos: -3.54896e+08 muA
** NormalTransistorPmos: -3.54897e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.9799e+08 muA
** DiodeTransistorPmos: -3.93389e+07 muA


** Expected Voltages: 
** ibias: 1.12801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.24501  V
** out: 2.5  V
** outFirstStage: 4.24901  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.22601  V
** innerStageBias: 0.503001  V
** innerTransistorStack1Load2: 0.613001  V
** innerTransistorStack2Load2: 0.612001  V
** sourceGCC1: 4.51301  V
** sourceGCC2: 4.51301  V
** sourceTransconductance: 1.86601  V
** innerStageBias: 0.573001  V
** innerTransconductance: 4.78201  V


.END