** Name: two_stage_single_output_op_amp_60_5

.MACRO two_stage_single_output_op_amp_60_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=16e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=187e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=17e-6
mMainBias5 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=2e-6 W=14e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=121e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=288e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=75e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=26e-6
mMainBias13 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mMainBias14 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=117e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=187e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=78e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=78e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=121e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=17e-6
mMainBias20 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=14e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=288e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=73e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_60_5

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 5.22201 mW
** Area: 7579 (mu_m)^2
** Transit frequency: 4.30001 MHz
** Transit frequency with error factor: 4.30033 MHz
** Slew rate: 4.62155 V/mu_s
** Phase margin: 69.328°
** CMRR: 143 dB
** VoutMax: 3.23001 V
** VoutMin: 0.540001 V
** VcmMax: 3.21001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.04801e+06 muA
** NormalTransistorNmos: 4.47341e+07 muA
** NormalTransistorNmos: 2.09031e+07 muA
** NormalTransistorNmos: 3.16171e+07 muA
** NormalTransistorNmos: 2.09031e+07 muA
** NormalTransistorNmos: 3.16171e+07 muA
** NormalTransistorPmos: -2.09039e+07 muA
** NormalTransistorPmos: -2.09039e+07 muA
** DiodeTransistorPmos: -2.09039e+07 muA
** NormalTransistorPmos: -2.14309e+07 muA
** DiodeTransistorPmos: -2.14319e+07 muA
** NormalTransistorPmos: -1.07149e+07 muA
** NormalTransistorPmos: -1.07149e+07 muA
** NormalTransistorNmos: 9.23286e+08 muA
** NormalTransistorPmos: -9.23285e+08 muA
** DiodeTransistorPmos: -9.23286e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.04899e+06 muA
** NormalTransistorPmos: -3.04999e+06 muA
** DiodeTransistorPmos: -4.47349e+07 muA
** NormalTransistorPmos: -4.47359e+07 muA


** Expected Voltages: 
** ibias: 1.15201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.947001  V
** outInputVoltageBiasXXpXX1: 3.38201  V
** outInputVoltageBiasXXpXX2: 2.67001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19101  V
** outSourceVoltageBiasXXpXX2: 3.83501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.25901  V
** out1: 3.51601  V
** sourceGCC1: 0.528001  V
** sourceGCC2: 0.528001  V
** sourceTransconductance: 3.23901  V
** inner: 4.19101  V
** inner: 3.83001  V


.END