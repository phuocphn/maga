** Name: two_stage_single_output_op_amp_94_12

.MACRO two_stage_single_output_op_amp_94_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=30e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=62e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=565e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=12e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=52e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=111e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=149e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=149e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=62e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=565e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=111e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=37e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=600e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=516e-6
mTelescopicFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=52e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=568e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mTelescopicFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=80e-6
mMainBias21 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=76e-6
mMainBias22 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.5e-12
.EOM two_stage_single_output_op_amp_94_12

** Expected Performance Values: 
** Gain: 184 dB
** Power consumption: 13.8411 mW
** Area: 14929 (mu_m)^2
** Transit frequency: 7.70001 MHz
** Transit frequency with error factor: 7.70018 MHz
** Slew rate: 8.80045 V/mu_s
** Phase margin: 60.7336°
** CMRR: 140 dB
** VoutMax: 4.10001 V
** VoutMin: 1 V
** VcmMax: 3.79001 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 1.22841e+07 muA
** NormalTransistorNmos: 2.01787e+08 muA
** NormalTransistorPmos: -2.30728e+08 muA
** NormalTransistorPmos: -3.01739e+07 muA
** NormalTransistorNmos: 7.09471e+07 muA
** NormalTransistorNmos: 7.09471e+07 muA
** DiodeTransistorPmos: -7.09479e+07 muA
** NormalTransistorPmos: -7.09479e+07 muA
** NormalTransistorPmos: -7.09479e+07 muA
** NormalTransistorNmos: 1.72069e+08 muA
** NormalTransistorNmos: 7.09481e+07 muA
** NormalTransistorNmos: 7.09481e+07 muA
** NormalTransistorNmos: 2.14127e+09 muA
** DiodeTransistorNmos: 2.14127e+09 muA
** NormalTransistorPmos: -2.14126e+09 muA
** NormalTransistorPmos: -2.14126e+09 muA
** DiodeTransistorNmos: 2.30729e+08 muA
** NormalTransistorNmos: 2.30729e+08 muA
** DiodeTransistorNmos: 3.01731e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.22849e+07 muA
** DiodeTransistorPmos: -2.01786e+08 muA


** Expected Voltages: 
** ibias: 0.571001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.97901  V
** outInputVoltageBiasXXnXX1: 1.40601  V
** outSourceVoltageBiasXXnXX1: 0.703001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 3.61101  V
** outVoltageBiasXXpXX1: 3.53401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 4.32001  V
** out1: 3.75601  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.54301  V
** inner: 0.703001  V


.END