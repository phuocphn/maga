** Name: two_stage_single_output_op_amp_11_10

.MACRO two_stage_single_output_op_amp_11_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mSimpleFirstStageLoad2 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=208e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=299e-6
mSecondStage1StageBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
mSimpleFirstStageTransconductor5 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=55e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=53e-6
mMainBias7 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=165e-6
mSecondStage1StageBias8 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=574e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=55e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=299e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=350e-6
mSecondStage1Transconductor12 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=208e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.5e-12
.EOM two_stage_single_output_op_amp_11_10

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 7.88401 mW
** Area: 6635 (mu_m)^2
** Transit frequency: 5.98201 MHz
** Transit frequency with error factor: 5.97912 MHz
** Slew rate: 5.63796 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** negPSRR: 112 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 0.260001 V
** VcmMax: 3.90001 V
** VcmMin: 0.820001 V


** Expected Currents: 
** NormalTransistorNmos: 3.24909e+08 muA
** DiodeTransistorPmos: -5.23789e+07 muA
** DiodeTransistorPmos: -5.23799e+07 muA
** NormalTransistorPmos: -5.23789e+07 muA
** NormalTransistorPmos: -5.23799e+07 muA
** NormalTransistorNmos: 1.04756e+08 muA
** NormalTransistorNmos: 5.23781e+07 muA
** NormalTransistorNmos: 5.23781e+07 muA
** NormalTransistorNmos: 1.13719e+09 muA
** NormalTransistorPmos: -1.13718e+09 muA
** NormalTransistorPmos: -1.13719e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.24908e+08 muA


** Expected Voltages: 
** ibias: 0.670001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.01101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.49401  V
** innerSourceLoad1: 4.26401  V
** innerTransistorStack2Load1: 4.26301  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.57501  V


.END