** Name: two_stage_single_output_op_amp_36_11

.MACRO two_stage_single_output_op_amp_36_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=9e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=286e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=29e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad5 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=16e-6
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=299e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
mSimpleFirstStageTransconductor9 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=29e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=510e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=286e-6
mMainBias13 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=143e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=528e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=537e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=557e-6
mSecondStage1Transconductor19 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=595e-6
mSimpleFirstStageLoad20 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=16e-6
mMainBias21 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=324e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_36_11

** Expected Performance Values: 
** Gain: 148 dB
** Power consumption: 6.76601 mW
** Area: 10968 (mu_m)^2
** Transit frequency: 3.41401 MHz
** Transit frequency with error factor: 3.41291 MHz
** Slew rate: 3.50013 V/mu_s
** Phase margin: 75.6305°
** CMRR: 108 dB
** negPSRR: 118 dB
** posPSRR: 104 dB
** VoutMax: 4.46001 V
** VoutMin: 0.710001 V
** VcmMax: 3.96001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 1.43114e+08 muA
** NormalTransistorNmos: 5.27977e+08 muA
** NormalTransistorPmos: -1.5341e+08 muA
** DiodeTransistorPmos: -7.88799e+06 muA
** DiodeTransistorPmos: -7.88899e+06 muA
** NormalTransistorPmos: -7.88799e+06 muA
** NormalTransistorPmos: -7.88899e+06 muA
** NormalTransistorNmos: 1.57751e+07 muA
** DiodeTransistorNmos: 1.57741e+07 muA
** NormalTransistorNmos: 7.88701e+06 muA
** NormalTransistorNmos: 7.88701e+06 muA
** NormalTransistorNmos: 5.02823e+08 muA
** NormalTransistorNmos: 5.02822e+08 muA
** NormalTransistorPmos: -5.02822e+08 muA
** NormalTransistorPmos: -5.02823e+08 muA
** DiodeTransistorNmos: 1.53411e+08 muA
** NormalTransistorNmos: 1.53411e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.43113e+08 muA
** DiodeTransistorPmos: -5.27976e+08 muA


** Expected Voltages: 
** ibias: 1.125  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.07101  V
** out: 2.5  V
** outFirstStage: 4.11701  V
** outInputVoltageBiasXXnXX1: 1.13001  V
** outSourceVoltageBiasXXnXX1: 0.565001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.55301  V
** innerSourceLoad1: 4.28301  V
** innerTransistorStack2Load1: 4.28301  V
** sourceTransconductance: 1.93201  V
** innerStageBias: 0.570001  V
** innerTransconductance: 4.46701  V
** inner: 0.565001  V


.END