** Name: one_stage_single_output_op_amp54

.MACRO one_stage_single_output_op_amp54 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=12e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=5e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=130e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=42e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=42e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=153e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=153e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=97e-6
mFoldedCascodeFirstStageLoad11 out inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=130e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=432e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=121e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=121e-6
mMainBias15 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=57e-6
mMainBias16 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mFoldedCascodeFirstStageLoad17 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=432e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp54

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 1.89301 mW
** Area: 5908 (mu_m)^2
** Transit frequency: 5.14801 MHz
** Transit frequency with error factor: 5.1482 MHz
** Slew rate: 4.35702 V/mu_s
** Phase margin: 83.6519°
** CMRR: 148 dB
** VoutMax: 3.93001 V
** VoutMin: 0.360001 V
** VcmMax: 5.05001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorPmos: -6.36669e+07 muA
** NormalTransistorPmos: -2.12929e+07 muA
** NormalTransistorPmos: -8.77249e+07 muA
** NormalTransistorPmos: -1.36851e+08 muA
** NormalTransistorPmos: -8.77249e+07 muA
** NormalTransistorPmos: -1.36851e+08 muA
** NormalTransistorNmos: 8.77241e+07 muA
** NormalTransistorNmos: 8.77231e+07 muA
** NormalTransistorNmos: 8.77241e+07 muA
** NormalTransistorNmos: 8.77231e+07 muA
** NormalTransistorNmos: 9.82511e+07 muA
** NormalTransistorNmos: 4.91261e+07 muA
** NormalTransistorNmos: 4.91261e+07 muA
** DiodeTransistorNmos: 6.36661e+07 muA
** DiodeTransistorNmos: 2.12921e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.04301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.962001  V
** inputVoltageBiasXXnXX2: 0.559001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.08201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.562001  V
** innerTransistorStack1Load2: 0.357001  V
** innerTransistorStack2Load2: 0.357001  V
** sourceGCC1: 3.75701  V
** sourceGCC2: 3.75701  V
** sourceTransconductance: 1.94401  V


.END