** Name: two_stage_single_output_op_amp_75_12

.MACRO two_stage_single_output_op_amp_75_12 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=190e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=9e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
mMainBias4 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=209e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=49e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=25e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYinnerStageBias inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=130e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=190e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=86e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=86e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=57e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=209e-6
mFoldedCascodeFirstStageLoad15 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=44e-6
mMainBias16 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=174e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=449e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=446e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=446e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=556e-6
mMainBias21 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=169e-6
mMainBias22 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=210e-6
mMainBias23 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=28e-6
mSecondStage1Transconductor24 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=600e-6
mFoldedCascodeFirstStageLoad25 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=449e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.5e-12
.EOM two_stage_single_output_op_amp_75_12

** Expected Performance Values: 
** Gain: 173 dB
** Power consumption: 5.80001 mW
** Area: 14893 (mu_m)^2
** Transit frequency: 3.21001 MHz
** Transit frequency with error factor: 3.20986 MHz
** Slew rate: 3.64994 V/mu_s
** Phase margin: 61.3065°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 1 V
** VcmMax: 5.25 V
** VcmMin: 1.46001 V


** Expected Currents: 
** NormalTransistorNmos: 8.30401e+07 muA
** NormalTransistorPmos: -3.41709e+07 muA
** NormalTransistorPmos: -4.28529e+07 muA
** NormalTransistorPmos: -5.64799e+06 muA
** NormalTransistorPmos: -6.07849e+07 muA
** NormalTransistorPmos: -9.17789e+07 muA
** NormalTransistorPmos: -6.07849e+07 muA
** NormalTransistorPmos: -9.17789e+07 muA
** DiodeTransistorNmos: 6.07841e+07 muA
** NormalTransistorNmos: 6.07841e+07 muA
** NormalTransistorNmos: 6.07841e+07 muA
** NormalTransistorNmos: 6.19851e+07 muA
** NormalTransistorNmos: 6.19841e+07 muA
** NormalTransistorNmos: 3.09931e+07 muA
** NormalTransistorNmos: 3.09931e+07 muA
** NormalTransistorNmos: 7.90698e+08 muA
** DiodeTransistorNmos: 7.90697e+08 muA
** NormalTransistorPmos: -7.90697e+08 muA
** NormalTransistorPmos: -7.90698e+08 muA
** DiodeTransistorNmos: 3.41701e+07 muA
** NormalTransistorNmos: 3.41691e+07 muA
** DiodeTransistorNmos: 4.28521e+07 muA
** DiodeTransistorNmos: 5.64701e+06 muA
** DiodeTransistorPmos: -8.30409e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.40601  V
** inputVoltageBiasXXnXX2: 1.06701  V
** inputVoltageBiasXXnXX3: 0.588001  V
** out: 2.5  V
** outFirstStage: 4.15401  V
** outSourceVoltageBiasXXnXX1: 0.703001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.383001  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.91001  V
** innerTransconductance: 4.71801  V
** inner: 0.701001  V


.END