** Name: two_stage_single_output_op_amp_119_11

.MACRO two_stage_single_output_op_amp_119_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=9e-6
mMainBias2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=145e-6
mTelescopicFirstStageLoad4 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=47e-6
mTelescopicFirstStageLoad5 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=26e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=33e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mTelescopicFirstStageLoad8 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=23e-6
mTelescopicFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=239e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=32e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=32e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mMainBias13 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=272e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=23e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=574e-6
mTelescopicFirstStageStageBias17 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=108e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=26e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=435e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad21 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=47e-6
mMainBias22 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=429e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.30001e-12
.EOM two_stage_single_output_op_amp_119_11

** Expected Performance Values: 
** Gain: 182 dB
** Power consumption: 7.13201 mW
** Area: 14792 (mu_m)^2
** Transit frequency: 2.53201 MHz
** Transit frequency with error factor: 2.53209 MHz
** Slew rate: 21.7435 V/mu_s
** Phase margin: 60.1606°
** CMRR: 132 dB
** VoutMax: 3.83001 V
** VoutMin: 0.790001 V
** VcmMax: 3.71001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 1.70131e+07 muA
** NormalTransistorNmos: 5.64078e+08 muA
** NormalTransistorPmos: -2.1875e+08 muA
** NormalTransistorNmos: 8.76201e+06 muA
** NormalTransistorNmos: 8.76201e+06 muA
** DiodeTransistorPmos: -8.76299e+06 muA
** DiodeTransistorPmos: -8.76399e+06 muA
** NormalTransistorPmos: -8.76299e+06 muA
** NormalTransistorPmos: -8.76399e+06 muA
** NormalTransistorNmos: 2.36272e+08 muA
** NormalTransistorNmos: 2.36271e+08 muA
** NormalTransistorNmos: 8.76101e+06 muA
** NormalTransistorNmos: 8.76101e+06 muA
** NormalTransistorNmos: 5.99102e+08 muA
** NormalTransistorNmos: 5.99101e+08 muA
** NormalTransistorPmos: -5.99101e+08 muA
** NormalTransistorPmos: -5.99102e+08 muA
** DiodeTransistorNmos: 2.18751e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.70139e+07 muA
** DiodeTransistorPmos: -5.64077e+08 muA


** Expected Voltages: 
** ibias: 1.125  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.92701  V
** out: 2.5  V
** outFirstStage: 3.59901  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX1: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerOutputLoad2: 3.45601  V
** innerStageBias: 0.492001  V
** innerTransistorStack1Load2: 4.19701  V
** innerTransistorStack2Load2: 4.19701  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.491001  V
** innerTransconductance: 2.83301  V


.END