** Name: two_stage_single_output_op_amp_55_3

.MACRO two_stage_single_output_op_amp_55_3 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=51e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=12e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=68e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=68e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=8e-6 W=213e-6
mMainBias10 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=367e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=318e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=51e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerOutputLoad2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=164e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=162e-6
mSecondStage1StageBias17 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=534e-6
mFoldedCascodeFirstStageLoad18 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=164e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_55_3

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 9.73701 mW
** Area: 8762 (mu_m)^2
** Transit frequency: 11.7661 MHz
** Transit frequency with error factor: 11.766 MHz
** Slew rate: 13.4394 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 3.28001 V
** VoutMin: 0.550001 V
** VcmMax: 4.66001 V
** VcmMin: 0.770001 V


** Expected Currents: 
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorPmos: -6.65799e+07 muA
** NormalTransistorPmos: -1.01533e+08 muA
** NormalTransistorPmos: -6.65799e+07 muA
** NormalTransistorPmos: -1.01533e+08 muA
** DiodeTransistorNmos: 6.65791e+07 muA
** NormalTransistorNmos: 6.65781e+07 muA
** NormalTransistorNmos: 6.65791e+07 muA
** DiodeTransistorNmos: 6.65781e+07 muA
** NormalTransistorNmos: 6.99111e+07 muA
** NormalTransistorNmos: 3.49551e+07 muA
** NormalTransistorNmos: 3.49551e+07 muA
** NormalTransistorNmos: 1.61246e+09 muA
** NormalTransistorPmos: -1.61245e+09 muA
** NormalTransistorPmos: -1.61245e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.21839e+08 muA
** DiodeTransistorPmos: -1.21839e+08 muA


** Expected Voltages: 
** ibias: 0.582001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.955001  V
** outSourceVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.16001  V
** innerSourceLoad2: 0.580001  V
** innerTransistorStack1Load2: 0.579001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.90401  V
** innerStageBias: 3.34601  V


.END