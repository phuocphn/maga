** Name: one_stage_single_output_op_amp121

.MACRO one_stage_single_output_op_amp121 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=6e-6
mMainBias2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=39e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=7e-6
mTelescopicFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=155e-6
mTelescopicFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=82e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=62e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=62e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
mTelescopicFirstStageLoad11 out outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=82e-6
mMainBias12 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=67e-6
mTelescopicFirstStageStageBias13 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=161e-6
mTelescopicFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=127e-6
mTelescopicFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=127e-6
mTelescopicFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=127e-6
mTelescopicFirstStageLoad17 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=127e-6
mMainBias18 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=8e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp121

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 1.22001 mW
** Area: 3126 (mu_m)^2
** Transit frequency: 4.16401 MHz
** Transit frequency with error factor: 4.16432 MHz
** Slew rate: 7.64378 V/mu_s
** Phase margin: 85.9437°
** CMRR: 148 dB
** VoutMax: 4.63001 V
** VoutMin: 0.600001 V
** VcmMax: 5.07001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 6.65721e+07 muA
** NormalTransistorNmos: 1.40111e+07 muA
** NormalTransistorPmos: -7.45969e+07 muA
** NormalTransistorNmos: 3.93621e+07 muA
** NormalTransistorNmos: 3.93621e+07 muA
** NormalTransistorPmos: -3.93629e+07 muA
** NormalTransistorPmos: -3.93639e+07 muA
** NormalTransistorPmos: -3.93629e+07 muA
** NormalTransistorPmos: -3.93639e+07 muA
** NormalTransistorNmos: 1.53324e+08 muA
** NormalTransistorNmos: 1.53323e+08 muA
** NormalTransistorNmos: 3.93631e+07 muA
** NormalTransistorNmos: 3.93631e+07 muA
** DiodeTransistorNmos: 7.45961e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -6.65729e+07 muA
** DiodeTransistorPmos: -1.40119e+07 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.87401  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 2.65801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.606001  V
** innerTransistorStack1Load2: 4.62401  V
** innerTransistorStack2Load2: 4.62401  V
** out1: 4.24901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END