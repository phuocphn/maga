** Name: two_stage_single_output_op_amp_61_4

.MACRO two_stage_single_output_op_amp_61_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=10e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=82e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=25e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=58e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=289e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=289e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=534e-6
mSecondStage1Transconductor10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=256e-6
mFoldedCascodeFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=58e-6
mMainBias12 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=33e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=243e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=82e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=30e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=30e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=3e-6 W=201e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=600e-6
mMainBias19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=164e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=600e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=103e-6
mMainBias22 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.4001e-12
.EOM two_stage_single_output_op_amp_61_4

** Expected Performance Values: 
** Gain: 180 dB
** Power consumption: 2.92501 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 3.14801 MHz
** Transit frequency with error factor: 3.14785 MHz
** Slew rate: 4.19953 V/mu_s
** Phase margin: 60.1606°
** CMRR: 136 dB
** VoutMax: 4.48001 V
** VoutMin: 0.330001 V
** VcmMax: 3.02001 V
** VcmMin: -0.369999 V


** Expected Currents: 
** NormalTransistorNmos: 1.35361e+07 muA
** NormalTransistorPmos: -6.67049e+07 muA
** NormalTransistorPmos: -4.02599e+06 muA
** NormalTransistorNmos: 6.90531e+07 muA
** NormalTransistorNmos: 1.18379e+08 muA
** NormalTransistorNmos: 6.90501e+07 muA
** NormalTransistorNmos: 1.18374e+08 muA
** DiodeTransistorPmos: -6.90519e+07 muA
** NormalTransistorPmos: -6.90509e+07 muA
** NormalTransistorPmos: -6.90519e+07 muA
** NormalTransistorPmos: -9.86489e+07 muA
** NormalTransistorPmos: -9.86499e+07 muA
** NormalTransistorPmos: -4.93239e+07 muA
** NormalTransistorPmos: -4.93239e+07 muA
** NormalTransistorNmos: 2.44045e+08 muA
** NormalTransistorNmos: 2.44044e+08 muA
** NormalTransistorPmos: -2.44042e+08 muA
** NormalTransistorPmos: -2.44041e+08 muA
** DiodeTransistorNmos: 6.67041e+07 muA
** DiodeTransistorNmos: 4.02501e+06 muA
** DiodeTransistorPmos: -1.35369e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.968001  V
** out: 2.5  V
** outFirstStage: 0.585001  V
** outVoltageBiasXXnXX2: 0.601001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.53601  V
** innerTransistorStack2Load2: 4.58401  V
** out1: 4.22001  V
** sourceGCC1: 0.396001  V
** sourceGCC2: 0.396001  V
** sourceTransconductance: 3.36601  V
** innerStageBias: 4.51101  V
** innerTransconductance: 0.413001  V


.END