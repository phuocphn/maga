** Name: two_stage_single_output_op_amp_176_1

.MACRO two_stage_single_output_op_amp_176_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=11e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=61e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=61e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=62e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mSimpleFirstStageLoad7 FirstStageYout1 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=446e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad9 outFirstStage ibias sourceNmos sourceNmos nmos4 L=9e-6 W=446e-6
mMainBias10 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=73e-6
mMainBias11 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=207e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=61e-6
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=247e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=600e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
mSecondStage1StageBias16 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=184e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=61e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=247e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.5e-12
.EOM two_stage_single_output_op_amp_176_1

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 12.3701 mW
** Area: 14499 (mu_m)^2
** Transit frequency: 13.6721 MHz
** Transit frequency with error factor: 13.6414 MHz
** Slew rate: 32.9679 V/mu_s
** Phase margin: 60.1606°
** CMRR: 75 dB
** VoutMax: 4.34001 V
** VoutMin: 0.170001 V
** VcmMax: 3 V
** VcmMin: -0.25 V


** Expected Currents: 
** NormalTransistorNmos: 6.58441e+07 muA
** NormalTransistorNmos: 1.87565e+08 muA
** DiodeTransistorPmos: -7.40939e+07 muA
** NormalTransistorPmos: -7.40949e+07 muA
** NormalTransistorPmos: -7.40939e+07 muA
** DiodeTransistorPmos: -7.40949e+07 muA
** NormalTransistorNmos: 3.99138e+08 muA
** NormalTransistorNmos: 3.99138e+08 muA
** NormalTransistorPmos: -6.50087e+08 muA
** DiodeTransistorPmos: -6.50087e+08 muA
** NormalTransistorPmos: -3.25043e+08 muA
** NormalTransistorPmos: -3.25043e+08 muA
** NormalTransistorNmos: 1.4124e+09 muA
** NormalTransistorPmos: -1.41239e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.58449e+07 muA
** NormalTransistorPmos: -6.58459e+07 muA
** DiodeTransistorPmos: -1.87564e+08 muA


** Expected Voltages: 
** ibias: 0.715001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.571001  V
** outInputVoltageBiasXXpXX1: 3.38201  V
** outSourceVoltageBiasXXpXX1: 4.19101  V
** outVoltageBiasXXpXX2: 3.77801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.85101  V
** innerTransistorStack1Load1: 3.84901  V
** out1: 3.02501  V
** sourceTransconductance: 3.44601  V
** inner: 4.18901  V


.END