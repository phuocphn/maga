** Name: symmetrical_op_amp56

.MACRO symmetrical_op_amp56 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=10e-6 W=14e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=45e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=45e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=56e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=1e-6 W=56e-6
mSymmetricalFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=85e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=10e-6 W=20e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=10e-6 W=20e-6
mSymmetricalFirstStageStageBias12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=85e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias13 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=56e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias15 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=56e-6
mSymmetricalFirstStageTransconductor16 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=143e-6
mSecondStage1StageBias17 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=56e-6
mSymmetricalFirstStageTransconductor18 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=143e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp56

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 1.30101 mW
** Area: 2252 (mu_m)^2
** Transit frequency: 3.45301 MHz
** Transit frequency with error factor: 3.45281 MHz
** Slew rate: 4.85294 V/mu_s
** Phase margin: 82.506°
** CMRR: 144 dB
** negPSRR: 40 dB
** posPSRR: 42 dB
** VoutMax: 3.99001 V
** VoutMin: 0.690001 V
** VcmMax: 3.17001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorPmos: -5.63339e+07 muA
** DiodeTransistorNmos: 4.30891e+07 muA
** DiodeTransistorNmos: 4.30891e+07 muA
** NormalTransistorPmos: -8.61799e+07 muA
** DiodeTransistorPmos: -8.61789e+07 muA
** NormalTransistorPmos: -4.30899e+07 muA
** NormalTransistorPmos: -4.30899e+07 muA
** NormalTransistorNmos: 4.85691e+07 muA
** NormalTransistorNmos: 4.85681e+07 muA
** NormalTransistorPmos: -4.85699e+07 muA
** DiodeTransistorPmos: -4.85709e+07 muA
** DiodeTransistorPmos: -4.90599e+07 muA
** NormalTransistorPmos: -4.90609e+07 muA
** NormalTransistorNmos: 4.90591e+07 muA
** NormalTransistorNmos: 4.90581e+07 muA
** DiodeTransistorNmos: 5.63331e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39601  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 1.09101  V
** inSourceStageBiasComplementarySecondStage: 4.21501  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 3.43001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.28801  V
** innerTransconductance: 0.150001  V
** inner: 4.21501  V
** inner: 0.150001  V
** inner: 4.19601  V


.END