** Name: two_stage_single_output_op_amp_100_3

.MACRO two_stage_single_output_op_amp_100_3 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=96e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=36e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos4 L=1e-6 W=19e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=94e-6
mTelescopicFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=573e-6
mMainBias6 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=4e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=304e-6
mTelescopicFirstStageLoad9 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=96e-6
mMainBias10 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mMainBias11 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=34e-6
mTelescopicFirstStageLoad12 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=4e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=284e-6
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=284e-6
mSecondStage1StageBias15 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=94e-6
mMainBias17 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=1e-6 W=85e-6
mSecondStage1StageBias18 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=600e-6
mTelescopicFirstStageLoad19 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=4e-6
mTelescopicFirstStageStageBias20 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=573e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.2001e-12
.EOM two_stage_single_output_op_amp_100_3

** Expected Performance Values: 
** Gain: 109 dB
** Power consumption: 4.73201 mW
** Area: 11464 (mu_m)^2
** Transit frequency: 6.875 MHz
** Transit frequency with error factor: 6.87225 MHz
** Slew rate: 11.2046 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** VoutMax: 3.96001 V
** VoutMin: 0.150001 V
** VcmMax: 3.03001 V
** VcmMin: 1.85001 V


** Expected Currents: 
** NormalTransistorNmos: 3.31181e+07 muA
** NormalTransistorNmos: 8.20521e+07 muA
** NormalTransistorPmos: -8.61789e+07 muA
** NormalTransistorPmos: -6.11369e+07 muA
** NormalTransistorPmos: -6.11369e+07 muA
** DiodeTransistorNmos: 6.11361e+07 muA
** NormalTransistorNmos: 6.11361e+07 muA
** NormalTransistorPmos: -2.04325e+08 muA
** DiodeTransistorPmos: -2.04326e+08 muA
** NormalTransistorPmos: -6.11359e+07 muA
** NormalTransistorPmos: -6.11359e+07 muA
** NormalTransistorNmos: 6.02852e+08 muA
** NormalTransistorPmos: -6.02851e+08 muA
** NormalTransistorPmos: -6.02852e+08 muA
** DiodeTransistorNmos: 8.61781e+07 muA
** DiodeTransistorPmos: -3.31189e+07 muA
** NormalTransistorPmos: -3.31199e+07 muA
** DiodeTransistorPmos: -8.20529e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.46301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.573001  V
** out: 2.5  V
** outFirstStage: 0.558001  V
** outInputVoltageBiasXXpXX1: 3.18001  V
** outSourceVoltageBiasXXpXX1: 4.09101  V
** outSourceVoltageBiasXXpXX3: 4.19901  V
** outVoltageBiasXXpXX2: 0.514001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21901  V
** out1: 0.555001  V
** sourceGCC1: 2.93601  V
** sourceGCC2: 2.93601  V
** innerStageBias: 4.26301  V
** inner: 4.08701  V


.END