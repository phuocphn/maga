** Name: two_stage_single_output_op_amp_9_9

.MACRO two_stage_single_output_op_amp_9_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=17e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=140e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=10e-6 W=205e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=9e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=9e-6 W=28e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=140e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=9e-6
mMainBias11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mSimpleFirstStageLoad12 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=10e-6 W=205e-6
mMainBias13 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=73e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=367e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=10e-6 W=33e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_9_9

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 3.01101 mW
** Area: 8305 (mu_m)^2
** Transit frequency: 3.22901 MHz
** Transit frequency with error factor: 3.22626 MHz
** Slew rate: 3.65561 V/mu_s
** Phase margin: 61.8795°
** CMRR: 100 dB
** negPSRR: 96 dB
** posPSRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 1 V
** VcmMax: 4.32001 V
** VcmMin: 0.830001 V


** Expected Currents: 
** NormalTransistorNmos: 5.19701e+06 muA
** NormalTransistorPmos: -3.82229e+07 muA
** NormalTransistorPmos: -8.24799e+06 muA
** NormalTransistorPmos: -8.24799e+06 muA
** DiodeTransistorPmos: -8.24799e+06 muA
** NormalTransistorNmos: 1.64931e+07 muA
** NormalTransistorNmos: 8.24701e+06 muA
** NormalTransistorNmos: 8.24701e+06 muA
** NormalTransistorNmos: 5.32328e+08 muA
** DiodeTransistorNmos: 5.32327e+08 muA
** NormalTransistorPmos: -5.32327e+08 muA
** DiodeTransistorNmos: 3.82221e+07 muA
** NormalTransistorNmos: 3.82211e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.19799e+06 muA


** Expected Voltages: 
** ibias: 0.654001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.40801  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.704001  V
** outVoltageBiasXXpXX0: 4.19401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.28601  V
** out1: 3.34901  V
** sourceTransconductance: 1.91401  V
** inner: 0.701001  V


.END