** Name: two_stage_single_output_op_amp_5_6

.MACRO two_stage_single_output_op_amp_5_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=28e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=232e-6
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=35e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=121e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=121e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=353e-6
mSecondStage1Transconductor10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=306e-6
mSimpleFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=35e-6
mMainBias12 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=81e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=55e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=560e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=28e-6
mMainBias16 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=460e-6
mSecondStage1StageBias17 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=232e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=55e-6
mMainBias19 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=44e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.10001e-12
.EOM two_stage_single_output_op_amp_5_6

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 5.33201 mW
** Area: 8133 (mu_m)^2
** Transit frequency: 17.0991 MHz
** Transit frequency with error factor: 17.0779 MHz
** Slew rate: 26.7187 V/mu_s
** Phase margin: 60.1606°
** CMRR: 101 dB
** negPSRR: 99 dB
** posPSRR: 224 dB
** VoutMax: 3.03001 V
** VoutMin: 0.380001 V
** VcmMax: 3.91001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 8.11461e+07 muA
** NormalTransistorPmos: -1.21129e+07 muA
** NormalTransistorPmos: -1.25078e+08 muA
** NormalTransistorNmos: 7.70861e+07 muA
** NormalTransistorNmos: 7.70851e+07 muA
** NormalTransistorNmos: 7.70861e+07 muA
** NormalTransistorNmos: 7.70851e+07 muA
** NormalTransistorPmos: -1.54173e+08 muA
** NormalTransistorPmos: -7.70869e+07 muA
** NormalTransistorPmos: -7.70869e+07 muA
** NormalTransistorNmos: 6.73969e+08 muA
** NormalTransistorNmos: 6.73968e+08 muA
** NormalTransistorPmos: -6.73968e+08 muA
** DiodeTransistorPmos: -6.73969e+08 muA
** DiodeTransistorNmos: 1.21121e+07 muA
** DiodeTransistorNmos: 1.25079e+08 muA
** DiodeTransistorPmos: -8.11469e+07 muA
** NormalTransistorPmos: -8.11479e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.782001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.47001  V
** outSourceVoltageBiasXXpXX1: 3.73501  V
** outVoltageBiasXXnXX0: 0.559001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.34301  V
** innerTransconductance: 0.150001  V
** inner: 3.72901  V


.END