** Name: two_stage_single_output_op_amp_134_3

.MACRO two_stage_single_output_op_amp_134_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=11e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=36e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=36e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=65e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=476e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=476e-6
mSimpleFirstStageLoad9 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=137e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=53e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=114e-6
mSimpleFirstStageLoad12 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=137e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=144e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=36e-6
mSimpleFirstStageTransconductor15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=31e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=86e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=577e-6
mSecondStage1StageBias18 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=471e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=36e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=31e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_134_3

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 5.84401 mW
** Area: 9178 (mu_m)^2
** Transit frequency: 4.15401 MHz
** Transit frequency with error factor: 4.14532 MHz
** Slew rate: 19.6756 V/mu_s
** Phase margin: 72.1927°
** CMRR: 90 dB
** VoutMax: 4.28001 V
** VoutMin: 0.360001 V
** VcmMax: 3.34001 V
** VcmMin: -0.129999 V


** Expected Currents: 
** NormalTransistorNmos: 2.53821e+07 muA
** NormalTransistorNmos: 6.90161e+07 muA
** DiodeTransistorPmos: -1.8276e+08 muA
** DiodeTransistorPmos: -1.8276e+08 muA
** NormalTransistorPmos: -1.8276e+08 muA
** NormalTransistorPmos: -1.8276e+08 muA
** NormalTransistorNmos: 2.27726e+08 muA
** NormalTransistorNmos: 2.27725e+08 muA
** NormalTransistorNmos: 2.27726e+08 muA
** NormalTransistorNmos: 2.27725e+08 muA
** NormalTransistorPmos: -8.99309e+07 muA
** NormalTransistorPmos: -4.49649e+07 muA
** NormalTransistorPmos: -4.49649e+07 muA
** NormalTransistorNmos: 6.08861e+08 muA
** NormalTransistorPmos: -6.0886e+08 muA
** NormalTransistorPmos: -6.08861e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.53829e+07 muA
** DiodeTransistorPmos: -6.90169e+07 muA


** Expected Voltages: 
** ibias: 1.16701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.762001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX2: 4.09301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.481001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.481001  V
** out1: 2.37201  V
** sourceTransconductance: 3.81401  V
** innerStageBias: 4.62901  V


.END