** Name: two_stage_single_output_op_amp_94_9

.MACRO two_stage_single_output_op_amp_94_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=599e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=5e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=127e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=70e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=35e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=35e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=599e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=70e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=6e-6 W=123e-6
mTelescopicFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=127e-6
mMainBias18 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=60e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=398e-6
mTelescopicFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=439e-6
mMainBias21 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.2001e-12
.EOM two_stage_single_output_op_amp_94_9

** Expected Performance Values: 
** Gain: 142 dB
** Power consumption: 14.9991 mW
** Area: 4512 (mu_m)^2
** Transit frequency: 11.4671 MHz
** Transit frequency with error factor: 11.4668 MHz
** Slew rate: 12.3358 V/mu_s
** Phase margin: 60.1606°
** CMRR: 154 dB
** VoutMax: 4.37001 V
** VoutMin: 0.870001 V
** VcmMax: 4.36001 V
** VcmMin: 0.850001 V


** Expected Currents: 
** NormalTransistorNmos: 7.54201e+06 muA
** NormalTransistorNmos: 7.47701e+06 muA
** NormalTransistorPmos: -4.55029e+07 muA
** NormalTransistorPmos: -1.88589e+07 muA
** NormalTransistorNmos: 6.66621e+07 muA
** NormalTransistorNmos: 6.66621e+07 muA
** DiodeTransistorPmos: -6.66629e+07 muA
** NormalTransistorPmos: -6.66629e+07 muA
** NormalTransistorPmos: -6.66629e+07 muA
** NormalTransistorNmos: 1.52182e+08 muA
** NormalTransistorNmos: 6.66621e+07 muA
** NormalTransistorNmos: 6.66621e+07 muA
** NormalTransistorNmos: 2.7772e+09 muA
** DiodeTransistorNmos: 2.77719e+09 muA
** NormalTransistorPmos: -2.77719e+09 muA
** DiodeTransistorNmos: 4.55021e+07 muA
** NormalTransistorNmos: 4.55011e+07 muA
** DiodeTransistorNmos: 1.88581e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.54299e+06 muA
** DiodeTransistorPmos: -7.47799e+06 muA


** Expected Voltages: 
** ibias: 0.702001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.27601  V
** out: 2.5  V
** outFirstStage: 3.80801  V
** outSourceVoltageBiasXXnXX1: 0.638001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 4.23001  V
** outVoltageBiasXXpXX1: 3.87301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 4.59601  V
** out1: 4.26401  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.638001  V


.END