** Name: symmetrical_op_amp189

.MACRO symmetrical_op_amp189 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=9e-6
mSecondStage1StageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=1e-6 W=20e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias5 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=68e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=48e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias8 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=53e-6
mSecondStage1StageBias10 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=1e-6 W=20e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=53e-6
mMainBias12 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=101e-6
mSymmetricalFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=47e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=47e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=67e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=67e-6
mSymmetricalFirstStageLoad17 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=83e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=120e-6
mSecondStage1Transconductor19 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=120e-6
mSymmetricalFirstStageLoad20 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=83e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp189

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 1.37201 mW
** Area: 3338 (mu_m)^2
** Transit frequency: 5.08201 MHz
** Transit frequency with error factor: 5.08179 MHz
** Slew rate: 4.83018 V/mu_s
** Phase margin: 71.0468°
** CMRR: 144 dB
** negPSRR: 118 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 0.740001 V
** VcmMax: 4.81001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00448e+08 muA
** NormalTransistorPmos: -3.36499e+07 muA
** NormalTransistorPmos: -3.36509e+07 muA
** NormalTransistorPmos: -3.36499e+07 muA
** NormalTransistorPmos: -3.36509e+07 muA
** NormalTransistorNmos: 6.72971e+07 muA
** NormalTransistorNmos: 6.72961e+07 muA
** NormalTransistorNmos: 3.36491e+07 muA
** NormalTransistorNmos: 3.36491e+07 muA
** NormalTransistorNmos: 4.83751e+07 muA
** DiodeTransistorNmos: 4.83741e+07 muA
** NormalTransistorPmos: -4.83759e+07 muA
** NormalTransistorPmos: -4.8375e+07 muA
** DiodeTransistorNmos: 4.83751e+07 muA
** NormalTransistorNmos: 4.83741e+07 muA
** NormalTransistorPmos: -4.83759e+07 muA
** NormalTransistorPmos: -4.8375e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.00447e+08 muA


** Expected Voltages: 
** ibias: 1.125  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 0.574001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 1.14801  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.538001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.40001  V
** inner: 0.574001  V
** inner: 4.40001  V


.END