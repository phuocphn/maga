** Name: two_stage_single_output_op_amp_122_7

.MACRO two_stage_single_output_op_amp_122_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=275e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=294e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=115e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=43e-6
mTelescopicFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=17e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=24e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=24e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=275e-6
mMainBias11 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=162e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=17e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=25e-6
mTelescopicFirstStageStageBias15 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=294e-6
mTelescopicFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=81e-6
mTelescopicFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=81e-6
mTelescopicFirstStageLoad18 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=60e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=490e-6
mTelescopicFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=60e-6
mMainBias21 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=302e-6
mMainBias22 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=302e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_122_7

** Expected Performance Values: 
** Gain: 148 dB
** Power consumption: 2.84101 mW
** Area: 11665 (mu_m)^2
** Transit frequency: 3.06301 MHz
** Transit frequency with error factor: 3.06333 MHz
** Slew rate: 6.48961 V/mu_s
** Phase margin: 62.4525°
** CMRR: 133 dB
** VoutMax: 4.81001 V
** VoutMin: 0.220001 V
** VcmMax: 5.09001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 2.51571e+07 muA
** NormalTransistorNmos: 1.19891e+07 muA
** NormalTransistorPmos: -1.74591e+08 muA
** NormalTransistorPmos: -1.73591e+08 muA
** NormalTransistorNmos: 6.53001e+06 muA
** NormalTransistorNmos: 6.53001e+06 muA
** NormalTransistorPmos: -6.53099e+06 muA
** NormalTransistorPmos: -6.53199e+06 muA
** NormalTransistorPmos: -6.53099e+06 muA
** NormalTransistorPmos: -6.53199e+06 muA
** NormalTransistorNmos: 1.86655e+08 muA
** DiodeTransistorNmos: 1.86655e+08 muA
** NormalTransistorNmos: 6.53101e+06 muA
** NormalTransistorNmos: 6.53101e+06 muA
** NormalTransistorNmos: 1.5984e+08 muA
** NormalTransistorPmos: -1.59839e+08 muA
** DiodeTransistorNmos: 1.74592e+08 muA
** NormalTransistorNmos: 1.74592e+08 muA
** DiodeTransistorNmos: 1.73592e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.51579e+07 muA
** DiodeTransistorPmos: -1.19899e+07 muA


** Expected Voltages: 
** ibias: 0.622001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.70701  V
** out: 2.5  V
** outFirstStage: 4.24401  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 3.99501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.42701  V
** innerTransistorStack2Load2: 4.42701  V
** out1: 4.27101  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.555001  V


.END