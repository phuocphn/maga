** Name: two_stage_single_output_op_amp_96_9

.MACRO two_stage_single_output_op_amp_96_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=10e-6 W=40e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=422e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=50e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=45e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=59e-6
mTelescopicFirstStageLoad7 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=12e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=9e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=9e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=422e-6
mTelescopicFirstStageLoad12 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=12e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=62e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=592e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=10e-6 W=423e-6
mTelescopicFirstStageLoad16 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=48e-6
mTelescopicFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=63e-6
mTelescopicFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=48e-6
mMainBias21 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=14e-6
mMainBias22 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=278e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_96_9

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 3.42301 mW
** Area: 14942 (mu_m)^2
** Transit frequency: 2.68401 MHz
** Transit frequency with error factor: 2.68448 MHz
** Slew rate: 16.3271 V/mu_s
** Phase margin: 62.4525°
** CMRR: 136 dB
** VoutMax: 4.40001 V
** VoutMin: 0.700001 V
** VcmMax: 5.08001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorNmos: 1.51951e+07 muA
** NormalTransistorNmos: 1.4698e+08 muA
** NormalTransistorPmos: -4.81099e+06 muA
** NormalTransistorPmos: -9.42899e+07 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorPmos: -5.71499e+06 muA
** NormalTransistorPmos: -5.71599e+06 muA
** NormalTransistorPmos: -5.71499e+06 muA
** NormalTransistorPmos: -5.71599e+06 muA
** NormalTransistorNmos: 1.05717e+08 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 4.01877e+08 muA
** DiodeTransistorNmos: 4.01877e+08 muA
** NormalTransistorPmos: -4.01876e+08 muA
** DiodeTransistorNmos: 4.81001e+06 muA
** NormalTransistorNmos: 4.80901e+06 muA
** DiodeTransistorNmos: 9.42891e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.51959e+07 muA
** DiodeTransistorPmos: -1.46979e+08 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.83601  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 4.19701  V
** outVoltageBiasXXpXX1: 3.69301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.25701  V
** innerTransistorStack1Load2: 4.42001  V
** innerTransistorStack2Load2: 4.42001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.554001  V


.END