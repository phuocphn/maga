** Name: two_stage_single_output_op_amp_31_7

.MACRO two_stage_single_output_op_amp_31_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=106e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=43e-6
mSimpleFirstStageStageBias5 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=30e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=16e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=33e-6
mSecondStage1StageBias8 out ibias sourceNmos sourceNmos nmos4 L=6e-6 W=597e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=16e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=60e-6
mSimpleFirstStageLoad11 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=106e-6
mMainBias12 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=24e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=42e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=51e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_31_7

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 2.61901 mW
** Area: 6198 (mu_m)^2
** Transit frequency: 2.68501 MHz
** Transit frequency with error factor: 2.68168 MHz
** Slew rate: 4.74736 V/mu_s
** Phase margin: 60.7336°
** CMRR: 102 dB
** negPSRR: 92 dB
** posPSRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 0.220001 V
** VcmMax: 4.5 V
** VcmMin: 1.49001 V


** Expected Currents: 
** NormalTransistorNmos: 4.26211e+07 muA
** NormalTransistorPmos: -2.33519e+07 muA
** NormalTransistorPmos: -1.07269e+07 muA
** NormalTransistorPmos: -1.07269e+07 muA
** DiodeTransistorPmos: -1.07269e+07 muA
** NormalTransistorNmos: 2.14511e+07 muA
** NormalTransistorNmos: 2.14501e+07 muA
** NormalTransistorNmos: 1.07261e+07 muA
** NormalTransistorNmos: 1.07261e+07 muA
** NormalTransistorNmos: 4.26443e+08 muA
** NormalTransistorPmos: -4.26442e+08 muA
** DiodeTransistorNmos: 2.33511e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.26219e+07 muA


** Expected Voltages: 
** ibias: 0.629001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.804001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 3.81601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.224001  V
** innerTransistorStack2Load1: 4.28601  V
** out1: 3.53501  V
** sourceTransconductance: 1.81301  V


.END