** Name: two_stage_single_output_op_amp_62_9

.MACRO two_stage_single_output_op_amp_62_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=11e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=31e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=599e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=102e-6
mMainBias6 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=119e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=307e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=29e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=16e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mSecondStage1StageBias13 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=599e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=16e-6
mMainBias15 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=102e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=32e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=32e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=307e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=119e-6
mMainBias21 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=249e-6
mMainBias22 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=365e-6
mSecondStage1Transconductor23 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=476e-6
mFoldedCascodeFirstStageLoad24 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=126e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_62_9

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 6.86901 mW
** Area: 14927 (mu_m)^2
** Transit frequency: 4.29401 MHz
** Transit frequency with error factor: 4.2935 MHz
** Slew rate: 4.04369 V/mu_s
** Phase margin: 73.3387°
** CMRR: 139 dB
** VoutMax: 4.36001 V
** VoutMin: 0.700001 V
** VcmMax: 3.29001 V
** VcmMin: -0.209999 V


** Expected Currents: 
** NormalTransistorNmos: 9.81481e+07 muA
** NormalTransistorPmos: -2.09519e+07 muA
** NormalTransistorPmos: -3.09779e+07 muA
** NormalTransistorNmos: 1.83551e+07 muA
** NormalTransistorNmos: 3.14671e+07 muA
** NormalTransistorNmos: 1.83521e+07 muA
** NormalTransistorNmos: 3.14621e+07 muA
** DiodeTransistorPmos: -1.83539e+07 muA
** NormalTransistorPmos: -1.83529e+07 muA
** NormalTransistorPmos: -1.83539e+07 muA
** NormalTransistorPmos: -2.62229e+07 muA
** DiodeTransistorPmos: -2.62219e+07 muA
** NormalTransistorPmos: -1.31109e+07 muA
** NormalTransistorPmos: -1.31109e+07 muA
** NormalTransistorNmos: 1.14088e+09 muA
** DiodeTransistorNmos: 1.14088e+09 muA
** NormalTransistorPmos: -1.14087e+09 muA
** DiodeTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** DiodeTransistorNmos: 3.09771e+07 muA
** DiodeTransistorNmos: 3.09781e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -9.81489e+07 muA


** Expected Voltages: 
** ibias: 3.50701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11001  V
** inputVoltageBiasXXnXX2: 1.31401  V
** out: 2.5  V
** outFirstStage: 3.79901  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.756001  V
** outSourceVoltageBiasXXpXX1: 4.25401  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.40601  V
** out1: 4.18901  V
** sourceGCC1: 0.744001  V
** sourceGCC2: 0.744001  V
** sourceTransconductance: 3.27801  V
** inner: 0.555001  V
** inner: 4.25201  V


.END