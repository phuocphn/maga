** Name: two_stage_single_output_op_amp_67_2

.MACRO two_stage_single_output_op_amp_67_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=65e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=26e-6
mFoldedCascodeFirstStageLoad4 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerOutputLoad2 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=31e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=161e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=161e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=285e-6
mSecondStage1Transconductor11 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=266e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=31e-6
mMainBias13 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=53e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=307e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=499e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=499e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=600e-6
mMainBias19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=410e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=149e-6
mSecondStage1StageBias21 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=26e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.7001e-12
.EOM two_stage_single_output_op_amp_67_2

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 8.55601 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 5.19101 MHz
** Transit frequency with error factor: 5.19121 MHz
** Slew rate: 8.65195 V/mu_s
** Phase margin: 60.1606°
** CMRR: 120 dB
** VoutMax: 4.69001 V
** VoutMin: 0.360001 V
** VcmMax: 3.03001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -3.44177e+08 muA
** NormalTransistorPmos: -1.23801e+08 muA
** NormalTransistorNmos: 1.79252e+08 muA
** NormalTransistorNmos: 3.0729e+08 muA
** NormalTransistorNmos: 1.79248e+08 muA
** NormalTransistorNmos: 3.07284e+08 muA
** DiodeTransistorPmos: -1.7925e+08 muA
** NormalTransistorPmos: -1.79248e+08 muA
** NormalTransistorPmos: -1.79247e+08 muA
** DiodeTransistorPmos: -1.79248e+08 muA
** NormalTransistorPmos: -2.56074e+08 muA
** NormalTransistorPmos: -2.56075e+08 muA
** NormalTransistorPmos: -1.28036e+08 muA
** NormalTransistorPmos: -1.28036e+08 muA
** NormalTransistorNmos: 5.07053e+08 muA
** NormalTransistorNmos: 5.07052e+08 muA
** NormalTransistorPmos: -5.07052e+08 muA
** DiodeTransistorNmos: 3.44178e+08 muA
** DiodeTransistorNmos: 1.23802e+08 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.01601  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.611001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 2.62401  V
** innerStageBias: 4.40401  V
** innerTransistorStack1Load2: 3.80701  V
** innerTransistorStack2Load2: 3.81201  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.44201  V
** innerTransconductance: 0.461001  V


.END