** Name: two_stage_single_output_op_amp_10_11

.MACRO two_stage_single_output_op_amp_10_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=9e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=15e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=269e-6
mMainBias4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=103e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=29e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=254e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=287e-6
mMainBias9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=49e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=7e-6 W=415e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=29e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=354e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=269e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=587e-6
mSecondStage1Transconductor15 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad16 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=69e-6
mMainBias17 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=90e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11e-12
.EOM two_stage_single_output_op_amp_10_11

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 5.50201 mW
** Area: 11926 (mu_m)^2
** Transit frequency: 5.33601 MHz
** Transit frequency with error factor: 5.32258 MHz
** Slew rate: 10.222 V/mu_s
** Phase margin: 60.1606°
** CMRR: 95 dB
** negPSRR: 132 dB
** posPSRR: 93 dB
** VoutMax: 4.65001 V
** VoutMin: 0.510001 V
** VcmMax: 4.34001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorNmos: 5.35191e+07 muA
** NormalTransistorNmos: 3.93243e+08 muA
** NormalTransistorPmos: -4.59849e+07 muA
** DiodeTransistorPmos: -1.3923e+08 muA
** NormalTransistorPmos: -1.3923e+08 muA
** NormalTransistorPmos: -1.3923e+08 muA
** NormalTransistorNmos: 2.7846e+08 muA
** NormalTransistorNmos: 1.39231e+08 muA
** NormalTransistorNmos: 1.39231e+08 muA
** NormalTransistorNmos: 3.19144e+08 muA
** NormalTransistorNmos: 3.19143e+08 muA
** NormalTransistorPmos: -3.19143e+08 muA
** NormalTransistorPmos: -3.19144e+08 muA
** DiodeTransistorNmos: 4.59841e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.35199e+07 muA
** DiodeTransistorPmos: -3.93242e+08 muA


** Expected Voltages: 
** ibias: 0.660001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.92701  V
** out: 2.5  V
** outFirstStage: 4.26201  V
** outVoltageBiasXXnXX1: 0.911001  V
** outVoltageBiasXXpXX1: 3.69801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.26501  V
** innerTransistorStack2Load1: 4.59701  V
** sourceTransconductance: 1.34501  V
** innerStageBias: 0.255001  V
** innerTransconductance: 4.43401  V


.END