** Name: two_stage_single_output_op_amp_43_9

.MACRO two_stage_single_output_op_amp_43_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=4e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=12e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=395e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=43e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=8e-6 W=157e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=59e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=27e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=27e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=395e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=59e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=17e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=8e-6 W=439e-6
mMainBias16 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=60e-6
mMainBias17 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=97e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=375e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=43e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_43_9

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 2.49501 mW
** Area: 12757 (mu_m)^2
** Transit frequency: 2.65501 MHz
** Transit frequency with error factor: 2.645 MHz
** Slew rate: 6.21246 V/mu_s
** Phase margin: 60.1606°
** CMRR: 86 dB
** VoutMax: 4.36001 V
** VoutMin: 0.770001 V
** VcmMax: 3.90001 V
** VcmMin: -0.289999 V


** Expected Currents: 
** NormalTransistorPmos: -3.86599e+06 muA
** NormalTransistorPmos: -6.15599e+06 muA
** NormalTransistorNmos: 2.80941e+07 muA
** NormalTransistorNmos: 4.21401e+07 muA
** NormalTransistorNmos: 2.80941e+07 muA
** NormalTransistorNmos: 4.21401e+07 muA
** DiodeTransistorPmos: -2.80949e+07 muA
** NormalTransistorPmos: -2.80949e+07 muA
** NormalTransistorPmos: -2.80949e+07 muA
** NormalTransistorPmos: -1.40469e+07 muA
** NormalTransistorPmos: -1.40469e+07 muA
** NormalTransistorNmos: 3.84647e+08 muA
** DiodeTransistorNmos: 3.84646e+08 muA
** NormalTransistorPmos: -3.84646e+08 muA
** DiodeTransistorNmos: 3.86501e+06 muA
** NormalTransistorNmos: 3.86401e+06 muA
** DiodeTransistorNmos: 6.15501e+06 muA
** DiodeTransistorNmos: 6.15601e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.18001  V
** inputVoltageBiasXXnXX2: 1.23601  V
** out: 2.5  V
** outFirstStage: 3.79901  V
** outSourceVoltageBiasXXnXX1: 0.590001  V
** outSourceVoltageBiasXXnXX2: 0.676001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.82901  V
** sourceGCC1: 0.681001  V
** sourceGCC2: 0.681001  V
** sourceTransconductance: 3.43501  V
** inner: 0.590001  V


.END