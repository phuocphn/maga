** Name: two_stage_single_output_op_amp_53_9

.MACRO two_stage_single_output_op_amp_53_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=59e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=6e-6 W=32e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=17e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=116e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=31e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=59e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=29e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=63e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=17e-6
mSecondStage1StageBias13 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=116e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=32e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=79e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
mMainBias18 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=108e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=591e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=79e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.90001e-12
.EOM two_stage_single_output_op_amp_53_9

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 5.04201 mW
** Area: 8381 (mu_m)^2
** Transit frequency: 3.35501 MHz
** Transit frequency with error factor: 3.35462 MHz
** Slew rate: 3.5927 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 4.25 V
** VoutMin: 1.63001 V
** VcmMax: 5.17001 V
** VcmMin: 0.840001 V


** Expected Currents: 
** NormalTransistorPmos: -1.09497e+08 muA
** NormalTransistorPmos: -2.12909e+07 muA
** NormalTransistorPmos: -3.20839e+07 muA
** NormalTransistorPmos: -5.37349e+07 muA
** NormalTransistorPmos: -3.20839e+07 muA
** NormalTransistorPmos: -5.37349e+07 muA
** DiodeTransistorNmos: 3.20831e+07 muA
** DiodeTransistorNmos: 3.20821e+07 muA
** NormalTransistorNmos: 3.20831e+07 muA
** NormalTransistorNmos: 3.20821e+07 muA
** NormalTransistorNmos: 4.32991e+07 muA
** NormalTransistorNmos: 2.16501e+07 muA
** NormalTransistorNmos: 2.16501e+07 muA
** NormalTransistorNmos: 7.50083e+08 muA
** DiodeTransistorNmos: 7.50082e+08 muA
** NormalTransistorPmos: -7.50082e+08 muA
** DiodeTransistorNmos: 1.09498e+08 muA
** NormalTransistorNmos: 1.09497e+08 muA
** DiodeTransistorNmos: 2.12901e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.04001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 1.02001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.606001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.601001  V
** innerTransistorStack2Load2: 0.600001  V
** out1: 1.27201  V
** sourceGCC1: 4.11201  V
** sourceGCC2: 4.11201  V
** sourceTransconductance: 1.86401  V
** inner: 1.01601  V


.END