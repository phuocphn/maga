** Name: two_stage_single_output_op_amp_152_7

.MACRO two_stage_single_output_op_amp_152_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=7e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=28e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=149e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=21e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=355e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=7e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=21e-6
mMainBias12 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=18e-6
mSimpleFirstStageLoad13 FirstStageYinnerOutputLoad1 outInputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=14e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=148e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=148e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=347e-6
mSimpleFirstStageLoad17 outFirstStage outInputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=14e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_152_7

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 5.12701 mW
** Area: 4410 (mu_m)^2
** Transit frequency: 4.32101 MHz
** Transit frequency with error factor: 4.31875 MHz
** Slew rate: 4.07258 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** VoutMax: 4.25 V
** VoutMin: 0.300001 V
** VcmMax: 4.45001 V
** VcmMin: 0.850001 V


** Expected Currents: 
** NormalTransistorNmos: 4.52531e+07 muA
** DiodeTransistorNmos: 3.46511e+07 muA
** NormalTransistorNmos: 3.46521e+07 muA
** NormalTransistorNmos: 3.46511e+07 muA
** DiodeTransistorNmos: 3.46521e+07 muA
** NormalTransistorPmos: -4.46519e+07 muA
** NormalTransistorPmos: -4.46529e+07 muA
** NormalTransistorPmos: -4.46519e+07 muA
** NormalTransistorPmos: -4.46529e+07 muA
** NormalTransistorNmos: 1.99991e+07 muA
** NormalTransistorNmos: 1.00001e+07 muA
** NormalTransistorNmos: 1.00001e+07 muA
** NormalTransistorNmos: 8.80808e+08 muA
** NormalTransistorPmos: -8.80807e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.52539e+07 muA
** DiodeTransistorPmos: -4.52549e+07 muA


** Expected Voltages: 
** ibias: 0.702001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXpXX1: 3.12301  V
** outSourceVoltageBiasXXpXX1: 4.21001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerTransistorStack1Load1: 1.04801  V
** innerTransistorStack1Load2: 4.41601  V
** innerTransistorStack2Load1: 1.04801  V
** innerTransistorStack2Load2: 4.41601  V
** sourceTransconductance: 1.94501  V


.END