** Name: two_stage_single_output_op_amp_168_1

.MACRO two_stage_single_output_op_amp_168_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=12e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=83e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=63e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=149e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=383e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=14e-6
mSimpleFirstStageLoad7 FirstStageYout1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=213e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=409e-6
mSimpleFirstStageLoad9 outFirstStage ibias sourceNmos sourceNmos nmos4 L=7e-6 W=213e-6
mMainBias10 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=43e-6
mMainBias11 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=19e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=83e-6
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=84e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=383e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=149e-6
mSecondStage1StageBias16 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=346e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=63e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=84e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.5e-12
.EOM two_stage_single_output_op_amp_168_1

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 4.00701 mW
** Area: 14986 (mu_m)^2
** Transit frequency: 4.44701 MHz
** Transit frequency with error factor: 4.43687 MHz
** Slew rate: 4.83766 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 0.150001 V
** VcmMax: 3.14001 V
** VcmMin: -0.299999 V


** Expected Currents: 
** NormalTransistorNmos: 3.53411e+07 muA
** NormalTransistorNmos: 1.57931e+07 muA
** DiodeTransistorPmos: -1.3006e+08 muA
** DiodeTransistorPmos: -1.30061e+08 muA
** NormalTransistorPmos: -1.3006e+08 muA
** NormalTransistorPmos: -1.30061e+08 muA
** NormalTransistorNmos: 1.75063e+08 muA
** NormalTransistorNmos: 1.75063e+08 muA
** NormalTransistorPmos: -9.00049e+07 muA
** DiodeTransistorPmos: -9.00059e+07 muA
** NormalTransistorPmos: -4.50019e+07 muA
** NormalTransistorPmos: -4.50019e+07 muA
** NormalTransistorNmos: 3.90227e+08 muA
** NormalTransistorPmos: -3.90226e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.53419e+07 muA
** NormalTransistorPmos: -3.53429e+07 muA
** DiodeTransistorPmos: -1.57939e+07 muA


** Expected Voltages: 
** ibias: 0.667001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.30801  V
** outSourceVoltageBiasXXpXX1: 4.15401  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.92101  V
** innerTransistorStack2Load1: 3.91601  V
** out1: 2.76601  V
** sourceTransconductance: 3.23701  V
** inner: 4.15301  V


.END