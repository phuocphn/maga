** Name: one_stage_single_output_op_amp102

.MACRO one_stage_single_output_op_amp102 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
mMainBias3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=22e-6
mTelescopicFirstStageStageBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=503e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=7e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
mTelescopicFirstStageLoad7 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=36e-6
mMainBias8 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=41e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=92e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=71e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=71e-6
mMainBias12 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mMainBias13 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mTelescopicFirstStageLoad14 out outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=92e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=503e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp102

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 1.29901 mW
** Area: 2856 (mu_m)^2
** Transit frequency: 2.78501 MHz
** Transit frequency with error factor: 2.78548 MHz
** Slew rate: 11.6007 V/mu_s
** Phase margin: 85.9437°
** CMRR: 133 dB
** VoutMax: 3.08001 V
** VoutMin: 0.860001 V
** VcmMax: 3 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorNmos: 3.85951e+07 muA
** NormalTransistorPmos: -7.39299e+06 muA
** NormalTransistorPmos: -9.69189e+07 muA
** NormalTransistorPmos: -9.69199e+07 muA
** NormalTransistorNmos: 9.69181e+07 muA
** NormalTransistorNmos: 9.69191e+07 muA
** DiodeTransistorNmos: 9.69181e+07 muA
** NormalTransistorPmos: -2.32432e+08 muA
** DiodeTransistorPmos: -2.32431e+08 muA
** NormalTransistorPmos: -9.69189e+07 muA
** NormalTransistorPmos: -9.69189e+07 muA
** DiodeTransistorNmos: 7.39301e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -3.85959e+07 muA


** Expected Voltages: 
** ibias: 3.55101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.702001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.27601  V
** outVoltageBiasXXpXX2: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.61401  V
** innerSourceLoad2: 0.680001  V
** out1: 1.26301  V
** sourceGCC1: 2.98501  V
** sourceGCC2: 2.98501  V
** inner: 4.27401  V


.END