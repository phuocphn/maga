** Name: symmetrical_op_amp195

.MACRO symmetrical_op_amp195 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=5e-6
mSecondStage1StageBias2 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=29e-6
mSymmetricalFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=22e-6
mMainBias4 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mSymmetricalFirstStageStageBias5 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=22e-6
mMainBias6 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mSymmetricalFirstStageTransconductor7 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=78e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias8 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=29e-6
mSecondStage1StageBias9 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos4 L=1e-6 W=22e-6
mSymmetricalFirstStageTransconductor10 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=78e-6
mMainBias11 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSymmetricalFirstStageLoad12 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=10e-6
mSymmetricalFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=10e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=25e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=25e-6
mSymmetricalFirstStageLoad16 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=107e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=267e-6
mSecondStage1Transconductor18 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=267e-6
mSymmetricalFirstStageLoad19 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=107e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp195

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 0.957001 mW
** Area: 3913 (mu_m)^2
** Transit frequency: 4.73501 MHz
** Transit frequency with error factor: 4.73475 MHz
** Slew rate: 5.3983 V/mu_s
** Phase margin: 81.3601°
** CMRR: 143 dB
** negPSRR: 116 dB
** posPSRR: 64 dB
** VoutMax: 4.25 V
** VoutMin: 0.970001 V
** VcmMax: 4.81001 V
** VcmMin: 1.52001 V


** Expected Currents: 
** NormalTransistorNmos: 3.00221e+07 muA
** NormalTransistorPmos: -2.15809e+07 muA
** NormalTransistorPmos: -2.15819e+07 muA
** NormalTransistorPmos: -2.15809e+07 muA
** NormalTransistorPmos: -2.15819e+07 muA
** NormalTransistorNmos: 4.31611e+07 muA
** DiodeTransistorNmos: 4.31621e+07 muA
** NormalTransistorNmos: 2.15801e+07 muA
** NormalTransistorNmos: 2.15801e+07 muA
** NormalTransistorNmos: 5.41511e+07 muA
** DiodeTransistorNmos: 5.41501e+07 muA
** NormalTransistorPmos: -5.41519e+07 muA
** NormalTransistorPmos: -5.41509e+07 muA
** NormalTransistorNmos: 5.41511e+07 muA
** NormalTransistorPmos: -5.41519e+07 muA
** NormalTransistorPmos: -5.41509e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.00229e+07 muA


** Expected Voltages: 
** ibias: 1.33801  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** inStageBiasComplementarySecondStage: 0.796001  V
** innerComplementarySecondStage: 1.37101  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.670001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.91401  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V
** inner: 0.666001  V


.END