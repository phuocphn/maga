** Name: two_stage_single_output_op_amp_144_12

.MACRO two_stage_single_output_op_amp_144_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=34e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=36e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=348e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=28e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=92e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=34e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=108e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=36e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=348e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=28e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=92e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=101e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=319e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=319e-6
mSimpleFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=532e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=545e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=532e-6
mMainBias22 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=200e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.5e-12
.EOM two_stage_single_output_op_amp_144_12

** Expected Performance Values: 
** Gain: 140 dB
** Power consumption: 11.0841 mW
** Area: 8006 (mu_m)^2
** Transit frequency: 7.48701 MHz
** Transit frequency with error factor: 7.48403 MHz
** Slew rate: 7.11555 V/mu_s
** Phase margin: 60.1606°
** CMRR: 108 dB
** VoutMax: 4.25 V
** VoutMin: 1.17001 V
** VcmMax: 4.96001 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 1.11687e+08 muA
** NormalTransistorNmos: 2.09481e+07 muA
** NormalTransistorPmos: -1.49727e+08 muA
** NormalTransistorNmos: 1.81365e+08 muA
** NormalTransistorNmos: 1.81366e+08 muA
** DiodeTransistorNmos: 1.81365e+08 muA
** NormalTransistorPmos: -2.40752e+08 muA
** NormalTransistorPmos: -2.40753e+08 muA
** NormalTransistorPmos: -2.40753e+08 muA
** NormalTransistorPmos: -2.40753e+08 muA
** NormalTransistorNmos: 1.18778e+08 muA
** NormalTransistorNmos: 5.93881e+07 muA
** NormalTransistorNmos: 5.93881e+07 muA
** NormalTransistorNmos: 1.44287e+09 muA
** DiodeTransistorNmos: 1.44287e+09 muA
** NormalTransistorPmos: -1.44286e+09 muA
** NormalTransistorPmos: -1.44286e+09 muA
** DiodeTransistorNmos: 1.49728e+08 muA
** NormalTransistorNmos: 1.49727e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.11686e+08 muA
** DiodeTransistorPmos: -2.09489e+07 muA


** Expected Voltages: 
** ibias: 0.567001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.05101  V
** outInputVoltageBiasXXnXX1: 1.57401  V
** outSourceVoltageBiasXXnXX1: 0.787001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.14601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack1Load2: 4.40901  V
** innerTransistorStack2Load2: 4.40901  V
** out1: 2.11601  V
** sourceTransconductance: 1.94301  V
** innerTransconductance: 4.61501  V
** inner: 0.784001  V


.END