** Name: one_stage_single_output_op_amp61

.MACRO one_stage_single_output_op_amp61 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=13e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=138e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=103e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=236e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=236e-6
mFoldedCascodeFirstStageLoad9 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=103e-6
mMainBias10 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=38e-6
mMainBias11 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=14e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=125e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=138e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=83e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=83e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=146e-6
mFoldedCascodeFirstStageLoad17 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=223e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp61

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 1.76601 mW
** Area: 3932 (mu_m)^2
** Transit frequency: 2.53201 MHz
** Transit frequency with error factor: 2.53185 MHz
** Slew rate: 5.12114 V/mu_s
** Phase margin: 88.8085°
** CMRR: 137 dB
** VoutMax: 4.57001 V
** VoutMin: 0.75 V
** VcmMax: 3.06001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.53531e+07 muA
** NormalTransistorNmos: 9.17701e+06 muA
** NormalTransistorNmos: 1.0279e+08 muA
** NormalTransistorNmos: 1.54342e+08 muA
** NormalTransistorNmos: 1.0279e+08 muA
** NormalTransistorNmos: 1.54342e+08 muA
** DiodeTransistorPmos: -1.02789e+08 muA
** NormalTransistorPmos: -1.02789e+08 muA
** NormalTransistorPmos: -1.02789e+08 muA
** NormalTransistorPmos: -1.03106e+08 muA
** NormalTransistorPmos: -1.03107e+08 muA
** NormalTransistorPmos: -5.15529e+07 muA
** NormalTransistorPmos: -5.15529e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.53539e+07 muA
** DiodeTransistorPmos: -9.17799e+06 muA


** Expected Voltages: 
** ibias: 1.12801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.22101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.53001  V
** innerTransistorStack2Load2: 4.47601  V
** out1: 4.23101  V
** sourceGCC1: 0.534001  V
** sourceGCC2: 0.534001  V
** sourceTransconductance: 3.38601  V


.END