** Name: two_stage_single_output_op_amp_46_4

.MACRO two_stage_single_output_op_amp_46_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=231e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=112e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=3e-6 W=544e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=11e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=193e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=240e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=240e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=490e-6
mSecondStage1Transconductor11 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=594e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=193e-6
mMainBias13 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=83e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=112e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=94e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=94e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=413e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
mMainBias19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=110e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=595e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=544e-6
mMainBias22 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=485e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.5e-12
.EOM two_stage_single_output_op_amp_46_4

** Expected Performance Values: 
** Gain: 169 dB
** Power consumption: 10.9501 mW
** Area: 14961 (mu_m)^2
** Transit frequency: 5.14001 MHz
** Transit frequency with error factor: 5.14012 MHz
** Slew rate: 15.5049 V/mu_s
** Phase margin: 60.1606°
** CMRR: 123 dB
** VoutMax: 4.45001 V
** VoutMin: 0.410001 V
** VcmMax: 3.37001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.59681e+08 muA
** NormalTransistorPmos: -9.97029e+07 muA
** NormalTransistorPmos: -4.39969e+08 muA
** NormalTransistorNmos: 2.67182e+08 muA
** NormalTransistorNmos: 4.58027e+08 muA
** NormalTransistorNmos: 2.67178e+08 muA
** NormalTransistorNmos: 4.58021e+08 muA
** DiodeTransistorPmos: -2.67179e+08 muA
** DiodeTransistorPmos: -2.67178e+08 muA
** NormalTransistorPmos: -2.67177e+08 muA
** NormalTransistorPmos: -2.67178e+08 muA
** NormalTransistorPmos: -3.81687e+08 muA
** NormalTransistorPmos: -1.90843e+08 muA
** NormalTransistorPmos: -1.90843e+08 muA
** NormalTransistorNmos: 5.54512e+08 muA
** NormalTransistorNmos: 5.54511e+08 muA
** NormalTransistorPmos: -5.54511e+08 muA
** NormalTransistorPmos: -5.5451e+08 muA
** DiodeTransistorNmos: 9.97021e+07 muA
** DiodeTransistorNmos: 4.3997e+08 muA
** DiodeTransistorPmos: -1.5968e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.01001  V
** out: 2.5  V
** outFirstStage: 0.605001  V
** outVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 3.80101  V
** innerTransistorStack2Load2: 3.79901  V
** out1: 2.94901  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.81401  V
** innerStageBias: 4.47801  V
** innerTransconductance: 0.394001  V


.END