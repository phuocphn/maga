** Name: symmetrical_op_amp186

.MACRO symmetrical_op_amp186 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=12e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mMainBias3 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=13e-6
mSymmetricalFirstStageStageBias5 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=32e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=12e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias8 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=10e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=28e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias10 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=5e-6 W=86e-6
mSecondStage1StageBias11 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=85e-6
mSymmetricalFirstStageTransconductor12 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=28e-6
mMainBias13 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=7e-6 W=37e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=10e-6
mSymmetricalFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=10e-6 W=21e-6
mSymmetricalFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=10e-6 W=21e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=10e-6 W=58e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=10e-6 W=58e-6
mMainBias19 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=53e-6
mSymmetricalFirstStageLoad20 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=66e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor21 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=186e-6
mSecondStage1Transconductor22 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=186e-6
mSymmetricalFirstStageLoad23 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=66e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp186

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 0.919001 mW
** Area: 4831 (mu_m)^2
** Transit frequency: 3.89501 MHz
** Transit frequency with error factor: 3.89549 MHz
** Slew rate: 3.74513 V/mu_s
** Phase margin: 60.7336°
** CMRR: 145 dB
** negPSRR: 147 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 0.630001 V
** VcmMax: 4.81001 V
** VcmMin: 1.59001 V


** Expected Currents: 
** NormalTransistorNmos: 8.21901e+06 muA
** NormalTransistorNmos: 3.04591e+07 muA
** NormalTransistorPmos: -3.32659e+07 muA
** NormalTransistorPmos: -1.33339e+07 muA
** NormalTransistorPmos: -1.33349e+07 muA
** NormalTransistorPmos: -1.33339e+07 muA
** NormalTransistorPmos: -1.33349e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 2.66641e+07 muA
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 3.75631e+07 muA
** NormalTransistorNmos: 3.75621e+07 muA
** NormalTransistorPmos: -3.75639e+07 muA
** NormalTransistorPmos: -3.75629e+07 muA
** NormalTransistorNmos: 3.75631e+07 muA
** NormalTransistorNmos: 3.75621e+07 muA
** NormalTransistorPmos: -3.75639e+07 muA
** NormalTransistorPmos: -3.75629e+07 muA
** DiodeTransistorNmos: 3.32651e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.21999e+06 muA
** DiodeTransistorPmos: -3.04599e+07 muA


** Expected Voltages: 
** ibias: 0.667001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 1.03501  V
** inSourceTransconductanceComplementarySecondStage: 3.83701  V
** innerComplementarySecondStage: 0.874001  V
** out: 2.5  V
** out1FirstStage: 3.83701  V
** out2FirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 4.01501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.266001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.469001  V
** innerTransconductance: 4.40001  V
** inner: 0.469001  V
** inner: 4.40001  V


.END