** Name: two_stage_single_output_op_amp_137_1

.MACRO two_stage_single_output_op_amp_137_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=33e-6
mSimpleFirstStageLoad2 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=20e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=42e-6
mSimpleFirstStageLoad5 FirstStageYinnerOutputLoad1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=192e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=535e-6
mSimpleFirstStageLoad7 outFirstStage outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=192e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=43e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=307e-6
mSecondStage1StageBias11 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=20e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=43e-6
mMainBias14 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=74e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.1001e-12
.EOM two_stage_single_output_op_amp_137_1

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 1.96201 mW
** Area: 10042 (mu_m)^2
** Transit frequency: 2.53601 MHz
** Transit frequency with error factor: 2.524 MHz
** Slew rate: 4.50459 V/mu_s
** Phase margin: 60.1606°
** CMRR: 79 dB
** VoutMax: 4.84001 V
** VoutMin: 0.150001 V
** VcmMax: 3.89001 V
** VcmMin: -0.319999 V


** Expected Currents: 
** NormalTransistorPmos: -1.77029e+07 muA
** DiodeTransistorPmos: -6.76889e+07 muA
** NormalTransistorPmos: -6.76889e+07 muA
** NormalTransistorPmos: -6.76889e+07 muA
** DiodeTransistorPmos: -6.76889e+07 muA
** NormalTransistorNmos: 1.04477e+08 muA
** NormalTransistorNmos: 1.04477e+08 muA
** NormalTransistorPmos: -7.35769e+07 muA
** NormalTransistorPmos: -3.67879e+07 muA
** NormalTransistorPmos: -3.67879e+07 muA
** NormalTransistorNmos: 1.45646e+08 muA
** NormalTransistorPmos: -1.45644e+08 muA
** DiodeTransistorNmos: 1.77021e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX1: 0.645001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerSourceLoad1: 3.68601  V
** innerTransistorStack1Load1: 3.68601  V
** sourceTransconductance: 3.44201  V


.END