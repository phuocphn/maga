** Name: two_stage_single_output_op_amp_54_11

.MACRO two_stage_single_output_op_amp_54_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=29e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=17e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=17e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=59e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=600e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=174e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=29e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=555e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=90e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=405e-6
mMainBias20 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=277e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=40e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_54_11

** Expected Performance Values: 
** Gain: 182 dB
** Power consumption: 2.19101 mW
** Area: 12004 (mu_m)^2
** Transit frequency: 2.68101 MHz
** Transit frequency with error factor: 2.68107 MHz
** Slew rate: 3.56455 V/mu_s
** Phase margin: 67.0361°
** CMRR: 140 dB
** VoutMax: 4.60001 V
** VoutMin: 0.360001 V
** VcmMax: 5.08001 V
** VcmMin: 0.770001 V


** Expected Currents: 
** NormalTransistorNmos: 1.52301e+08 muA
** NormalTransistorNmos: 2.46321e+07 muA
** NormalTransistorPmos: -3.57939e+07 muA
** NormalTransistorPmos: -1.61069e+07 muA
** NormalTransistorPmos: -2.41589e+07 muA
** NormalTransistorPmos: -1.61109e+07 muA
** NormalTransistorPmos: -2.41649e+07 muA
** NormalTransistorNmos: 1.61081e+07 muA
** NormalTransistorNmos: 1.61091e+07 muA
** NormalTransistorNmos: 1.61101e+07 muA
** NormalTransistorNmos: 1.61091e+07 muA
** NormalTransistorNmos: 1.61071e+07 muA
** NormalTransistorNmos: 8.05301e+06 muA
** NormalTransistorNmos: 8.05301e+06 muA
** NormalTransistorNmos: 1.6711e+08 muA
** NormalTransistorNmos: 1.67109e+08 muA
** NormalTransistorPmos: -1.67109e+08 muA
** NormalTransistorPmos: -1.6711e+08 muA
** DiodeTransistorNmos: 3.57931e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.523e+08 muA
** DiodeTransistorPmos: -2.46329e+07 muA


** Expected Voltages: 
** ibias: 0.556001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.05201  V
** out: 2.5  V
** outFirstStage: 4.22101  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.11201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.690001  V
** innerTransistorStack1Load2: 0.485001  V
** innerTransistorStack2Load2: 0.485001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.88301  V
** innerStageBias: 0.433001  V
** innerTransconductance: 4.43301  V


.END