** Name: two_stage_single_output_op_amp_58_9

.MACRO two_stage_single_output_op_amp_58_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=32e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=24e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=450e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=46e-6
mMainBias6 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=63e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=394e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=18e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=32e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=450e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=18e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=196e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=196e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=394e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=63e-6
mMainBias18 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=444e-6
mMainBias19 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=329e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=407e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=46e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.5e-12
.EOM two_stage_single_output_op_amp_58_9

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 6.58801 mW
** Area: 14421 (mu_m)^2
** Transit frequency: 4.54801 MHz
** Transit frequency with error factor: 4.54164 MHz
** Slew rate: 4.65899 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 0.730001 V
** VcmMax: 3.22001 V
** VcmMin: -0.369999 V


** Expected Currents: 
** NormalTransistorPmos: -7.12599e+07 muA
** NormalTransistorPmos: -5.20449e+07 muA
** NormalTransistorNmos: 4.43281e+07 muA
** NormalTransistorNmos: 7.59921e+07 muA
** NormalTransistorNmos: 4.43261e+07 muA
** NormalTransistorNmos: 7.59881e+07 muA
** DiodeTransistorPmos: -4.43269e+07 muA
** NormalTransistorPmos: -4.43269e+07 muA
** NormalTransistorPmos: -6.33259e+07 muA
** DiodeTransistorPmos: -6.33249e+07 muA
** NormalTransistorPmos: -3.16629e+07 muA
** NormalTransistorPmos: -3.16629e+07 muA
** NormalTransistorNmos: 1.02231e+09 muA
** DiodeTransistorNmos: 1.02231e+09 muA
** NormalTransistorPmos: -1.0223e+09 muA
** DiodeTransistorNmos: 7.12591e+07 muA
** NormalTransistorNmos: 7.12581e+07 muA
** DiodeTransistorNmos: 5.20441e+07 muA
** DiodeTransistorNmos: 5.20431e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.44801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.13601  V
** inputVoltageBiasXXnXX2: 1.16701  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.568001  V
** outSourceVoltageBiasXXnXX2: 0.602001  V
** outSourceVoltageBiasXXpXX1: 4.22501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.69901  V
** sourceGCC1: 0.591001  V
** sourceGCC2: 0.591001  V
** sourceTransconductance: 3.29601  V
** inner: 0.568001  V
** inner: 4.22201  V


.END