** Name: two_stage_single_output_op_amp_206_12

.MACRO two_stage_single_output_op_amp_206_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=70e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=70e-6
mMainBias3 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=8e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=54e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=56e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=372e-6
mMainBias7 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=60e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mSimpleFirstStageTransconductor9 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=12e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=70e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=56e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=54e-6
mMainBias13 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mMainBias14 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=30e-6
mSecondStage1StageBias15 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=372e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=70e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=12e-6
mMainBias18 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mSimpleFirstStageLoad19 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=312e-6
mSimpleFirstStageLoad20 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=521e-6
mSimpleFirstStageLoad21 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=521e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=514e-6
mSecondStage1Transconductor23 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=503e-6
mSimpleFirstStageLoad24 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=312e-6
mMainBias25 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=35e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.20001e-12
.EOM two_stage_single_output_op_amp_206_12

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 5.86701 mW
** Area: 14992 (mu_m)^2
** Transit frequency: 4.56801 MHz
** Transit frequency with error factor: 4.56624 MHz
** Slew rate: 4.30539 V/mu_s
** Phase margin: 60.1606°
** CMRR: 124 dB
** VoutMax: 4.33001 V
** VoutMin: 0.890001 V
** VcmMax: 4.67001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00151e+07 muA
** NormalTransistorNmos: 3.68131e+07 muA
** NormalTransistorPmos: -2.18489e+07 muA
** DiodeTransistorNmos: 3.07735e+08 muA
** NormalTransistorNmos: 3.07736e+08 muA
** NormalTransistorNmos: 3.07737e+08 muA
** DiodeTransistorNmos: 3.07736e+08 muA
** NormalTransistorPmos: -3.19162e+08 muA
** NormalTransistorPmos: -3.19163e+08 muA
** NormalTransistorPmos: -3.19164e+08 muA
** NormalTransistorPmos: -3.19163e+08 muA
** NormalTransistorNmos: 2.28551e+07 muA
** DiodeTransistorNmos: 2.28541e+07 muA
** NormalTransistorNmos: 1.14281e+07 muA
** NormalTransistorNmos: 1.14281e+07 muA
** NormalTransistorNmos: 4.56478e+08 muA
** DiodeTransistorNmos: 4.56479e+08 muA
** NormalTransistorPmos: -4.56477e+08 muA
** NormalTransistorPmos: -4.56478e+08 muA
** DiodeTransistorNmos: 2.18481e+07 muA
** NormalTransistorNmos: 2.18471e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.00159e+07 muA
** DiodeTransistorPmos: -3.68139e+07 muA


** Expected Voltages: 
** ibias: 1.29201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.17301  V
** out: 2.5  V
** outFirstStage: 4.21201  V
** outInputVoltageBiasXXnXX1: 1.24801  V
** outSourceVoltageBiasXXnXX1: 0.624001  V
** outSourceVoltageBiasXXnXX2: 0.647001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.12901  V
** innerTransistorStack1Load1: 1.13001  V
** innerTransistorStack1Load2: 4.72701  V
** innerTransistorStack2Load2: 4.72701  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.69901  V
** inner: 0.624001  V
** inner: 0.643001  V


.END