** Name: two_stage_single_output_op_amp_93_7

.MACRO two_stage_single_output_op_amp_93_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=9e-6
mTelescopicFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=6e-6 W=90e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=16e-6
mTelescopicFirstStageLoad5 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=22e-6
mTelescopicFirstStageTransconductor6 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=11e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=11e-6
mSecondStage1StageBias8 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad9 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=22e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mTelescopicFirstStageStageBias11 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=53e-6
mTelescopicFirstStageLoad12 FirstStageYout1 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=6e-6 W=90e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=382e-6
mTelescopicFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=31e-6
mMainBias15 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=42e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.2001e-12
.EOM two_stage_single_output_op_amp_93_7

** Expected Performance Values: 
** Gain: 133 dB
** Power consumption: 4.78901 mW
** Area: 4307 (mu_m)^2
** Transit frequency: 4.35201 MHz
** Transit frequency with error factor: 4.35222 MHz
** Slew rate: 7.42466 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 4.38001 V
** VoutMin: 0.180001 V
** VcmMax: 4.07001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorNmos: 1.28851e+07 muA
** NormalTransistorPmos: -3.39449e+07 muA
** NormalTransistorNmos: 2.09521e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorPmos: -2.09529e+07 muA
** NormalTransistorPmos: -2.09519e+07 muA
** DiodeTransistorPmos: -2.09529e+07 muA
** NormalTransistorNmos: 7.58451e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 8.59044e+08 muA
** NormalTransistorPmos: -8.59043e+08 muA
** DiodeTransistorNmos: 3.39441e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.28859e+07 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.81901  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 3.79601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 4.15601  V
** out1: 3.25501  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END