** Name: two_stage_single_output_op_amp_15_6

.MACRO two_stage_single_output_op_amp_15_6 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=119e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=16e-6
mSecondStage1StageBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=4e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=429e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mSecondStage1Transconductor9 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=153e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=119e-6
mMainBias11 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mSimpleFirstStageStageBias12 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=75e-6
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=491e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=38e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mMainBias16 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias17 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=429e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=491e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=68e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_15_6

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 6.70201 mW
** Area: 11177 (mu_m)^2
** Transit frequency: 16.1891 MHz
** Transit frequency with error factor: 16.1774 MHz
** Slew rate: 16.401 V/mu_s
** Phase margin: 71.6198°
** CMRR: 101 dB
** negPSRR: 93 dB
** posPSRR: 95 dB
** VoutMax: 3.09001 V
** VoutMin: 0.570001 V
** VcmMax: 3.14001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 1.08761e+07 muA
** NormalTransistorPmos: -1.01379e+07 muA
** NormalTransistorPmos: -6.89429e+07 muA
** DiodeTransistorNmos: 3.80201e+07 muA
** NormalTransistorNmos: 3.80201e+07 muA
** NormalTransistorPmos: -7.60409e+07 muA
** NormalTransistorPmos: -7.60399e+07 muA
** NormalTransistorPmos: -3.80209e+07 muA
** NormalTransistorPmos: -3.80209e+07 muA
** NormalTransistorNmos: 1.15432e+09 muA
** NormalTransistorNmos: 1.15432e+09 muA
** NormalTransistorPmos: -1.15431e+09 muA
** DiodeTransistorPmos: -1.15432e+09 muA
** DiodeTransistorNmos: 1.01371e+07 muA
** DiodeTransistorNmos: 6.89421e+07 muA
** DiodeTransistorPmos: -1.08769e+07 muA
** NormalTransistorPmos: -1.08779e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.578001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.52201  V
** outSourceVoltageBiasXXpXX1: 3.76101  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX1: 0.976001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.29501  V
** out1: 0.555001  V
** sourceTransconductance: 3.22501  V
** innerTransconductance: 0.150001  V
** inner: 3.75901  V


.END