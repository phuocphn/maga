** Name: two_stage_single_output_op_amp_178_5

.MACRO two_stage_single_output_op_amp_178_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=8e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=13e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=3e-6 W=13e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=257e-6
mMainBias6 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=2e-6 W=37e-6
mSimpleFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=253e-6
mSecondStage1StageBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=135e-6
mSimpleFirstStageLoad9 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=79e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=114e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=114e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=236e-6
mSimpleFirstStageLoad13 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=79e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=44e-6
mMainBias15 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=350e-6
mSimpleFirstStageTransconductor16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=113e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=3e-6 W=13e-6
mSimpleFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=253e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=257e-6
mMainBias20 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=37e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=135e-6
mSimpleFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=13e-6
mSimpleFirstStageTransconductor23 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=113e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_178_5

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 4.57001 mW
** Area: 12962 (mu_m)^2
** Transit frequency: 3.80201 MHz
** Transit frequency with error factor: 3.79956 MHz
** Slew rate: 4.51024 V/mu_s
** Phase margin: 69.9009°
** CMRR: 103 dB
** VoutMax: 3.01001 V
** VoutMin: 0.390001 V
** VcmMax: 3.35001 V
** VcmMin: -0.229999 V


** Expected Currents: 
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 1.66656e+08 muA
** DiodeTransistorPmos: -4.39979e+07 muA
** NormalTransistorPmos: -4.39979e+07 muA
** NormalTransistorPmos: -4.39979e+07 muA
** DiodeTransistorPmos: -4.39979e+07 muA
** NormalTransistorNmos: 5.42811e+07 muA
** NormalTransistorNmos: 5.42821e+07 muA
** NormalTransistorNmos: 5.42811e+07 muA
** NormalTransistorNmos: 5.42821e+07 muA
** NormalTransistorPmos: -2.05689e+07 muA
** DiodeTransistorPmos: -2.05699e+07 muA
** NormalTransistorPmos: -1.02839e+07 muA
** NormalTransistorPmos: -1.02839e+07 muA
** NormalTransistorNmos: 6.07884e+08 muA
** NormalTransistorPmos: -6.07883e+08 muA
** DiodeTransistorPmos: -6.07884e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.09519e+07 muA
** NormalTransistorPmos: -2.09529e+07 muA
** DiodeTransistorPmos: -1.66655e+08 muA
** NormalTransistorPmos: -1.66656e+08 muA


** Expected Voltages: 
** ibias: 1.20201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.797001  V
** outInputVoltageBiasXXpXX1: 3.54001  V
** outInputVoltageBiasXXpXX2: 2.44601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.27001  V
** outSourceVoltageBiasXXpXX2: 3.72301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.616001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.616001  V
** sourceTransconductance: 3.25201  V
** inner: 4.26901  V
** inner: 3.71701  V


.END