** Name: two_stage_single_output_op_amp_6_6

.MACRO two_stage_single_output_op_amp_6_6 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=50e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=6e-6 W=50e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
mSecondStage1StageBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=8e-6 W=150e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=179e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=464e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=6e-6 W=50e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=32e-6
mSecondStage1Transconductor10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=512e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=50e-6
mMainBias12 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=202e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=37e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=8e-6 W=488e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=179e-6
mMainBias16 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=106e-6
mMainBias17 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=333e-6
mSecondStage1StageBias18 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=464e-6
mSimpleFirstStageTransconductor19 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=37e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.40001e-12
.EOM two_stage_single_output_op_amp_6_6

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 2.16101 mW
** Area: 14292 (mu_m)^2
** Transit frequency: 3.53201 MHz
** Transit frequency with error factor: 3.52751 MHz
** Slew rate: 6.06843 V/mu_s
** Phase margin: 60.1606°
** CMRR: 101 dB
** negPSRR: 103 dB
** posPSRR: 216 dB
** VoutMax: 4.09001 V
** VoutMin: 0.460001 V
** VcmMax: 3.99001 V
** VcmMin: 0.550001 V


** Expected Currents: 
** NormalTransistorNmos: 9.69901e+07 muA
** NormalTransistorPmos: -7.15799e+06 muA
** NormalTransistorPmos: -2.20729e+07 muA
** DiodeTransistorNmos: 1.64761e+07 muA
** NormalTransistorNmos: 1.64751e+07 muA
** NormalTransistorNmos: 1.64761e+07 muA
** DiodeTransistorNmos: 1.64751e+07 muA
** NormalTransistorPmos: -3.29539e+07 muA
** NormalTransistorPmos: -1.64769e+07 muA
** NormalTransistorPmos: -1.64769e+07 muA
** NormalTransistorNmos: 2.53102e+08 muA
** NormalTransistorNmos: 2.53101e+08 muA
** NormalTransistorPmos: -2.53101e+08 muA
** DiodeTransistorPmos: -2.53102e+08 muA
** DiodeTransistorNmos: 7.15701e+06 muA
** DiodeTransistorNmos: 2.20721e+07 muA
** DiodeTransistorPmos: -9.69909e+07 muA
** NormalTransistorPmos: -9.69919e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.555001  V
** inputVoltageBiasXXnXX1: 0.864001  V
** out: 2.5  V
** outFirstStage: 0.711001  V
** outInputVoltageBiasXXpXX1: 3.52201  V
** outSourceVoltageBiasXXpXX1: 4.26101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 1.11601  V
** innerTransistorStack1Load1: 0.558001  V
** innerTransistorStack2Load1: 0.558001  V
** sourceTransconductance: 3.33701  V
** innerTransconductance: 0.306001  V
** inner: 4.26001  V


.END