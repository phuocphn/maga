** Name: two_stage_single_output_op_amp_196_7

.MACRO two_stage_single_output_op_amp_196_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=6e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=5e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=146e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=70e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=146e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=591e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=6e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=70e-6
mSimpleFirstStageLoad14 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=236e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=404e-6
mSimpleFirstStageLoad16 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=236e-6
mMainBias17 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias18 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.6001e-12
.EOM two_stage_single_output_op_amp_196_7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 14.9991 mW
** Area: 4633 (mu_m)^2
** Transit frequency: 7.18901 MHz
** Transit frequency with error factor: 7.18166 MHz
** Slew rate: 6.77585 V/mu_s
** Phase margin: 60.1606°
** CMRR: 84 dB
** VoutMax: 4.38001 V
** VoutMin: 0.400001 V
** VcmMax: 5.25 V
** VcmMin: 1.42001 V


** Expected Currents: 
** NormalTransistorPmos: -4.52999e+06 muA
** NormalTransistorPmos: -1.82389e+07 muA
** DiodeTransistorNmos: 4.23901e+07 muA
** DiodeTransistorNmos: 4.23891e+07 muA
** NormalTransistorNmos: 4.23901e+07 muA
** NormalTransistorNmos: 4.23891e+07 muA
** NormalTransistorPmos: -1.09052e+08 muA
** NormalTransistorPmos: -1.09052e+08 muA
** NormalTransistorNmos: 1.33324e+08 muA
** DiodeTransistorNmos: 1.33323e+08 muA
** NormalTransistorNmos: 6.66621e+07 muA
** NormalTransistorNmos: 6.66621e+07 muA
** NormalTransistorNmos: 2.73903e+09 muA
** NormalTransistorPmos: -2.73902e+09 muA
** DiodeTransistorNmos: 4.52901e+06 muA
** NormalTransistorNmos: 4.52801e+06 muA
** DiodeTransistorNmos: 1.82401e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.81701  V
** outInputVoltageBiasXXnXX1: 1.27401  V
** outSourceVoltageBiasXXnXX1: 0.637001  V
** outVoltageBiasXXnXX2: 0.809001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.11001  V
** innerTransistorStack2Load1: 1.10401  V
** out1: 2.15801  V
** sourceTransconductance: 1.94501  V
** inner: 0.637001  V


.END