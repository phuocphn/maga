** Name: two_stage_single_output_op_amp_63_2

.MACRO two_stage_single_output_op_amp_63_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=112e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=64e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mMainBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=177e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=470e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=470e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=535e-6
mMainBias11 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=191e-6
mSecondStage1Transconductor12 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=535e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=177e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=252e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=112e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=430e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=430e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=519e-6
mMainBias19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=145e-6
mSecondStage1StageBias20 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=64e-6
mMainBias22 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.2001e-12
.EOM two_stage_single_output_op_amp_63_2

** Expected Performance Values: 
** Gain: 131 dB
** Power consumption: 6.94701 mW
** Area: 14988 (mu_m)^2
** Transit frequency: 7.56901 MHz
** Transit frequency with error factor: 7.569 MHz
** Slew rate: 13.5186 V/mu_s
** Phase margin: 60.1606°
** CMRR: 123 dB
** VoutMax: 4.78001 V
** VoutMin: 0.300001 V
** VcmMax: 3.20001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorPmos: -1.22319e+08 muA
** NormalTransistorPmos: -1.84129e+07 muA
** NormalTransistorNmos: 1.93192e+08 muA
** NormalTransistorNmos: 2.98393e+08 muA
** NormalTransistorNmos: 1.93192e+08 muA
** NormalTransistorNmos: 2.98393e+08 muA
** DiodeTransistorPmos: -1.93191e+08 muA
** DiodeTransistorPmos: -1.93192e+08 muA
** NormalTransistorPmos: -1.93191e+08 muA
** NormalTransistorPmos: -1.93192e+08 muA
** NormalTransistorPmos: -2.104e+08 muA
** NormalTransistorPmos: -2.10401e+08 muA
** NormalTransistorPmos: -1.05199e+08 muA
** NormalTransistorPmos: -1.05199e+08 muA
** NormalTransistorNmos: 5.09989e+08 muA
** NormalTransistorNmos: 5.09988e+08 muA
** NormalTransistorPmos: -5.09987e+08 muA
** DiodeTransistorNmos: 1.2232e+08 muA
** DiodeTransistorNmos: 1.84121e+07 muA
** DiodeTransistorPmos: -1.21839e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.915001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40001  V
** innerTransistorStack1Load2: 3.89601  V
** innerTransistorStack2Load2: 3.89001  V
** out1: 2.61701  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.37301  V
** innerTransconductance: 0.360001  V


.END