** Name: two_stage_single_output_op_amp_167_5

.MACRO two_stage_single_output_op_amp_167_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=23e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=166e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=62e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=349e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=78e-6
mSimpleFirstStageLoad8 FirstStageYout1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mMainBias9 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=153e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=517e-6
mSimpleFirstStageLoad11 outFirstStage ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mMainBias12 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=380e-6
mSimpleFirstStageStageBias13 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=535e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=323e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=597e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
mSecondStage1StageBias18 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=349e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=23e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=323e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.2001e-12
.EOM two_stage_single_output_op_amp_167_5

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 9.13001 mW
** Area: 14135 (mu_m)^2
** Transit frequency: 12.2001 MHz
** Transit frequency with error factor: 12.1705 MHz
** Slew rate: 28.0332 V/mu_s
** Phase margin: 60.1606°
** CMRR: 70 dB
** VoutMax: 3.64001 V
** VoutMin: 0.150001 V
** VcmMax: 3.02001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorNmos: 1.79061e+08 muA
** NormalTransistorNmos: 7.23811e+07 muA
** DiodeTransistorPmos: -4.20989e+07 muA
** DiodeTransistorPmos: -4.20999e+07 muA
** NormalTransistorPmos: -4.20989e+07 muA
** NormalTransistorPmos: -4.20999e+07 muA
** NormalTransistorNmos: 2.86158e+08 muA
** NormalTransistorNmos: 2.86158e+08 muA
** NormalTransistorPmos: -4.88117e+08 muA
** NormalTransistorPmos: -4.88118e+08 muA
** NormalTransistorPmos: -2.44058e+08 muA
** NormalTransistorPmos: -2.44058e+08 muA
** NormalTransistorNmos: 9.92151e+08 muA
** NormalTransistorPmos: -9.9215e+08 muA
** DiodeTransistorPmos: -9.92151e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.7906e+08 muA
** NormalTransistorPmos: -1.79059e+08 muA
** DiodeTransistorPmos: -7.23819e+07 muA
** DiodeTransistorPmos: -7.23829e+07 muA


** Expected Voltages: 
** ibias: 0.572001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.48901  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.07201  V
** outSourceVoltageBiasXXpXX1: 4.03601  V
** outSourceVoltageBiasXXpXX2: 4.20901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.94901  V
** innerStageBias: 4.26601  V
** innerTransistorStack2Load1: 3.94701  V
** out1: 3.06401  V
** sourceTransconductance: 3.47401  V
** inner: 4.03701  V


.END