** Name: two_stage_single_output_op_amp_151_8

.MACRO two_stage_single_output_op_amp_151_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
mMainBias4 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=61e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=45e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=358e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=241e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=10e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=45e-6
mSimpleFirstStageLoad13 FirstStageYinnerOutputLoad1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=396e-6
mMainBias14 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=493e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=233e-6
mSimpleFirstStageLoad16 outFirstStage ibias sourcePmos sourcePmos pmos4 L=3e-6 W=396e-6
mMainBias17 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=452e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.9001e-12
.EOM two_stage_single_output_op_amp_151_8

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 7.44701 mW
** Area: 7430 (mu_m)^2
** Transit frequency: 3.78701 MHz
** Transit frequency with error factor: 3.77905 MHz
** Slew rate: 3.56898 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** VoutMax: 4.25 V
** VoutMin: 0.540001 V
** VcmMax: 5.24001 V
** VcmMin: 0.75 V


** Expected Currents: 
** NormalTransistorPmos: -7.45239e+07 muA
** NormalTransistorPmos: -8.13179e+07 muA
** DiodeTransistorNmos: 4.39611e+07 muA
** NormalTransistorNmos: 4.39621e+07 muA
** NormalTransistorNmos: 4.39631e+07 muA
** DiodeTransistorNmos: 4.39621e+07 muA
** NormalTransistorPmos: -6.53899e+07 muA
** NormalTransistorPmos: -6.53899e+07 muA
** NormalTransistorNmos: 4.28551e+07 muA
** NormalTransistorNmos: 2.14281e+07 muA
** NormalTransistorNmos: 2.14281e+07 muA
** NormalTransistorNmos: 1.18288e+09 muA
** NormalTransistorNmos: 1.18288e+09 muA
** NormalTransistorPmos: -1.18287e+09 muA
** DiodeTransistorNmos: 7.45231e+07 muA
** DiodeTransistorNmos: 8.13171e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.602001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 0.944001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.12901  V
** innerTransistorStack1Load1: 1.13001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.197001  V


.END