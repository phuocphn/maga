** Name: two_stage_single_output_op_amp_123_9

.MACRO two_stage_single_output_op_amp_123_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=10e-6 W=21e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=289e-6
mMainBias4 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=27e-6
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mTelescopicFirstStageLoad7 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=10e-6
mMainBias8 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=15e-6
mTelescopicFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=416e-6
mTelescopicFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=9e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=6e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=6e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=289e-6
mTelescopicFirstStageLoad16 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=9e-6
mTelescopicFirstStageStageBias17 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=105e-6
mTelescopicFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=340e-6
mTelescopicFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=10e-6
mMainBias21 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=75e-6
mMainBias22 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=535e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_123_9

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 3.20201 mW
** Area: 12995 (mu_m)^2
** Transit frequency: 2.69101 MHz
** Transit frequency with error factor: 2.69137 MHz
** Slew rate: 17.605 V/mu_s
** Phase margin: 60.7336°
** CMRR: 138 dB
** VoutMax: 4.10001 V
** VoutMin: 0.820001 V
** VcmMax: 3.70001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorNmos: 1.92301e+06 muA
** NormalTransistorPmos: -9.47499e+06 muA
** NormalTransistorPmos: -6.78889e+07 muA
** NormalTransistorNmos: 5.71501e+06 muA
** NormalTransistorNmos: 5.71501e+06 muA
** DiodeTransistorPmos: -5.71599e+06 muA
** NormalTransistorPmos: -5.71699e+06 muA
** NormalTransistorPmos: -5.71599e+06 muA
** DiodeTransistorPmos: -5.71699e+06 muA
** NormalTransistorNmos: 7.93151e+07 muA
** NormalTransistorNmos: 7.93141e+07 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.397e+08 muA
** DiodeTransistorNmos: 5.39699e+08 muA
** NormalTransistorPmos: -5.39699e+08 muA
** DiodeTransistorNmos: 9.47401e+06 muA
** NormalTransistorNmos: 9.47301e+06 muA
** DiodeTransistorNmos: 6.78881e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.92399e+06 muA


** Expected Voltages: 
** ibias: 1.19601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.26701  V
** out: 2.5  V
** outFirstStage: 3.53801  V
** outInputVoltageBiasXXnXX1: 1.23001  V
** outSourceVoltageBiasXXnXX1: 0.616001  V
** outSourceVoltageBiasXXnXX3: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.18201  V
** innerStageBias: 0.491001  V
** innerTransistorStack1Load2: 4.18101  V
** out1: 3.43901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.613001  V


.END