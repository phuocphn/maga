** Name: two_stage_single_output_op_amp_61_12

.MACRO two_stage_single_output_op_amp_61_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=11e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=514e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=9e-6 W=203e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=22e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=38e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=38e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=514e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=22e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=39e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=9e-6 W=329e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=120e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=120e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=13e-6
mSecondStage1Transconductor20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=523e-6
mMainBias21 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=9e-6 W=142e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=598e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=72e-6
mMainBias24 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=9e-6 W=387e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_61_12

** Expected Performance Values: 
** Gain: 177 dB
** Power consumption: 5.49401 mW
** Area: 14995 (mu_m)^2
** Transit frequency: 3.29501 MHz
** Transit frequency with error factor: 3.29547 MHz
** Slew rate: 3.5193 V/mu_s
** Phase margin: 79.0682°
** CMRR: 144 dB
** VoutMax: 4.25 V
** VoutMin: 0.700001 V
** VcmMax: 3.17001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.50101e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -6.98499e+06 muA
** NormalTransistorNmos: 1.59321e+07 muA
** NormalTransistorNmos: 2.41261e+07 muA
** NormalTransistorNmos: 1.59321e+07 muA
** NormalTransistorNmos: 2.41261e+07 muA
** DiodeTransistorPmos: -1.59329e+07 muA
** NormalTransistorPmos: -1.59329e+07 muA
** NormalTransistorPmos: -1.59329e+07 muA
** NormalTransistorPmos: -1.63909e+07 muA
** NormalTransistorPmos: -1.63919e+07 muA
** NormalTransistorPmos: -8.19499e+06 muA
** NormalTransistorPmos: -8.19499e+06 muA
** NormalTransistorNmos: 9.79444e+08 muA
** DiodeTransistorNmos: 9.79443e+08 muA
** NormalTransistorPmos: -9.79443e+08 muA
** NormalTransistorPmos: -9.79444e+08 muA
** DiodeTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** DiodeTransistorNmos: 6.98401e+06 muA
** DiodeTransistorNmos: 6.98401e+06 muA
** DiodeTransistorPmos: -2.50109e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.11001  V
** out: 2.5  V
** outFirstStage: 4.11201  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.62401  V
** innerTransistorStack2Load2: 4.40701  V
** out1: 4.21301  V
** sourceGCC1: 0.544001  V
** sourceGCC2: 0.544001  V
** sourceTransconductance: 3.23801  V
** innerTransconductance: 4.67601  V
** inner: 0.555001  V


.END