** Name: two_stage_single_output_op_amp_89_9

.MACRO two_stage_single_output_op_amp_89_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=22e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=575e-6
mMainBias4 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=63e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=5e-6
mTelescopicFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=16e-6
mTelescopicFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=48e-6
mTelescopicFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=48e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=575e-6
mTelescopicFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=16e-6
mMainBias13 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=11e-6
mTelescopicFirstStageLoad14 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=5e-6 W=127e-6
mTelescopicFirstStageTransconductor15 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=29e-6
mTelescopicFirstStageTransconductor16 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=29e-6
mMainBias17 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=350e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=368e-6
mTelescopicFirstStageLoad19 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=5e-6 W=127e-6
mMainBias20 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=121e-6
mMainBias21 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=14e-6
mTelescopicFirstStageStageBias22 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=5e-6 W=144e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.20001e-12
.EOM two_stage_single_output_op_amp_89_9

** Expected Performance Values: 
** Gain: 131 dB
** Power consumption: 11.6611 mW
** Area: 11031 (mu_m)^2
** Transit frequency: 2.54901 MHz
** Transit frequency with error factor: 2.54863 MHz
** Slew rate: 4.41183 V/mu_s
** Phase margin: 60.1606°
** CMRR: 150 dB
** VoutMax: 3.46001 V
** VoutMin: 1 V
** VcmMax: 3.98001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 2.71801e+06 muA
** NormalTransistorPmos: -2.24399e+06 muA
** NormalTransistorPmos: -1.91509e+07 muA
** NormalTransistorPmos: -5.53169e+07 muA
** NormalTransistorPmos: -1.02139e+07 muA
** NormalTransistorPmos: -1.02129e+07 muA
** NormalTransistorNmos: 1.02131e+07 muA
** NormalTransistorNmos: 1.02121e+07 muA
** NormalTransistorNmos: 1.02121e+07 muA
** NormalTransistorNmos: 1.02121e+07 muA
** NormalTransistorPmos: -2.31439e+07 muA
** NormalTransistorPmos: -1.02129e+07 muA
** NormalTransistorPmos: -1.02129e+07 muA
** NormalTransistorNmos: 2.21245e+09 muA
** DiodeTransistorNmos: 2.21245e+09 muA
** NormalTransistorPmos: -2.21244e+09 muA
** DiodeTransistorNmos: 2.24301e+06 muA
** DiodeTransistorNmos: 1.91501e+07 muA
** NormalTransistorNmos: 1.91491e+07 muA
** DiodeTransistorNmos: 5.53161e+07 muA
** DiodeTransistorPmos: -2.71899e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.22501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.705001  V
** out: 2.5  V
** outFirstStage: 2.89401  V
** outInputVoltageBiasXXnXX1: 1.41001  V
** outSourceVoltageBiasXXnXX1: 0.705001  V
** outVoltageBiasXXnXX0: 0.567001  V
** outVoltageBiasXXpXX1: 2.35001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.30601  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 3.06401  V
** sourceGCC2: 3.06401  V
** inner: 0.705001  V


.END