** Name: two_stage_single_output_op_amp_1_6

.MACRO two_stage_single_output_op_amp_1_6 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=119e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mSecondStage1StageBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=5e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=407e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=425e-6
mSecondStage1Transconductor8 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=302e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=119e-6
mMainBias10 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=15e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=28e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=600e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias14 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=19e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=163e-6
mSecondStage1StageBias16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=407e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=28e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_1_6

** Expected Performance Values: 
** Gain: 133 dB
** Power consumption: 5.18701 mW
** Area: 7212 (mu_m)^2
** Transit frequency: 13.6491 MHz
** Transit frequency with error factor: 13.6217 MHz
** Slew rate: 32.8233 V/mu_s
** Phase margin: 67.6091°
** CMRR: 93 dB
** negPSRR: 88 dB
** posPSRR: 93 dB
** VoutMax: 3.49001 V
** VoutMin: 0.460001 V
** VcmMax: 3.81001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 1.01371e+07 muA
** NormalTransistorPmos: -4.80299e+06 muA
** NormalTransistorPmos: -4.08439e+07 muA
** DiodeTransistorNmos: 7.60401e+07 muA
** NormalTransistorNmos: 7.60401e+07 muA
** NormalTransistorPmos: -1.5208e+08 muA
** NormalTransistorPmos: -7.60409e+07 muA
** NormalTransistorPmos: -7.60409e+07 muA
** NormalTransistorNmos: 8.09468e+08 muA
** NormalTransistorNmos: 8.09467e+08 muA
** NormalTransistorPmos: -8.09467e+08 muA
** DiodeTransistorPmos: -8.09468e+08 muA
** DiodeTransistorNmos: 4.80201e+06 muA
** DiodeTransistorNmos: 4.08431e+07 muA
** DiodeTransistorPmos: -1.01379e+07 muA
** NormalTransistorPmos: -1.01379e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.642001  V
** inputVoltageBiasXXnXX1: 0.862001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.92401  V
** outSourceVoltageBiasXXpXX1: 3.96201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceTransconductance: 3.45201  V
** innerTransconductance: 0.150001  V
** inner: 3.96201  V


.END