** Name: two_stage_single_output_op_amp_114_10

.MACRO two_stage_single_output_op_amp_114_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=25e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=209e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=99e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=48e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=453e-6
mSecondStage1StageBias7 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=11e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=11e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=11e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=25e-6
mMainBias12 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mMainBias13 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=243e-6
mSecondStage1StageBias14 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=508e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=11e-6
mTelescopicFirstStageStageBias16 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=209e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=493e-6
mSecondStage1Transconductor18 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=273e-6
mTelescopicFirstStageLoad19 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=48e-6
mMainBias20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=73e-6
mMainBias21 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=581e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_114_10

** Expected Performance Values: 
** Gain: 107 dB
** Power consumption: 5.45101 mW
** Area: 13580 (mu_m)^2
** Transit frequency: 4.92301 MHz
** Transit frequency with error factor: 4.91998 MHz
** Slew rate: 9.62345 V/mu_s
** Phase margin: 61.8795°
** CMRR: 82 dB
** VoutMax: 4.52001 V
** VoutMin: 0.170001 V
** VcmMax: 4.53001 V
** VcmMin: 1.56001 V


** Expected Currents: 
** NormalTransistorNmos: 2.8594e+08 muA
** NormalTransistorNmos: 1.15895e+08 muA
** NormalTransistorPmos: -4.66349e+07 muA
** NormalTransistorPmos: -3.73382e+08 muA
** NormalTransistorNmos: 1.04761e+07 muA
** NormalTransistorNmos: 1.04761e+07 muA
** DiodeTransistorPmos: -1.04769e+07 muA
** NormalTransistorPmos: -1.04769e+07 muA
** NormalTransistorNmos: 3.94334e+08 muA
** DiodeTransistorNmos: 3.94333e+08 muA
** NormalTransistorNmos: 1.04761e+07 muA
** NormalTransistorNmos: 1.04761e+07 muA
** NormalTransistorNmos: 2.37484e+08 muA
** NormalTransistorPmos: -2.37483e+08 muA
** NormalTransistorPmos: -2.37484e+08 muA
** DiodeTransistorNmos: 4.66341e+07 muA
** NormalTransistorNmos: 4.66331e+07 muA
** DiodeTransistorNmos: 3.73383e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.85939e+08 muA
** DiodeTransistorPmos: -1.15894e+08 muA


** Expected Voltages: 
** ibias: 0.572001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.10901  V
** inputVoltageBiasXXpXX1: 2.81801  V
** out: 2.5  V
** outFirstStage: 4.27101  V
** outInputVoltageBiasXXnXX1: 1.40601  V
** outSourceVoltageBiasXXnXX1: 0.703001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.27901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 3.69301  V
** inner: 0.703001  V


.END