** Name: symmetrical_op_amp97

.MACRO symmetrical_op_amp97 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mMainBias2 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=54e-6
mSecondStage1StageBias3 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=27e-6
mSymmetricalFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=27e-6
mSecondStage1Transconductor6 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=47e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor7 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=47e-6
mSymmetricalFirstStageLoad8 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=43e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=65e-6
mSecondStage1Transconductor10 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=65e-6
mSymmetricalFirstStageLoad11 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=43e-6
mSymmetricalFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=5e-6 W=552e-6
mSymmetricalFirstStageTransconductor13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=208e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias14 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias15 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=1e-6 W=161e-6
mSymmetricalFirstStageTransconductor16 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=208e-6
mMainBias17 out2FirstStage ibias sourcePmos sourcePmos pmos4 L=5e-6 W=95e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp97

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 1.60201 mW
** Area: 6414 (mu_m)^2
** Transit frequency: 7 MHz
** Transit frequency with error factor: 6.99961 MHz
** Slew rate: 8.92789 V/mu_s
** Phase margin: 79.6412°
** CMRR: 149 dB
** negPSRR: 46 dB
** posPSRR: 68 dB
** VoutMax: 3.55001 V
** VoutMin: 0.460001 V
** VcmMax: 4 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.78279e+07 muA
** NormalTransistorNmos: 5.17951e+07 muA
** NormalTransistorNmos: 5.17941e+07 muA
** NormalTransistorNmos: 5.17951e+07 muA
** NormalTransistorNmos: 5.17941e+07 muA
** NormalTransistorPmos: -1.03591e+08 muA
** NormalTransistorPmos: -5.17959e+07 muA
** NormalTransistorPmos: -5.17959e+07 muA
** NormalTransistorNmos: 8.95171e+07 muA
** NormalTransistorNmos: 8.95181e+07 muA
** NormalTransistorPmos: -8.95179e+07 muA
** DiodeTransistorPmos: -8.95189e+07 muA
** NormalTransistorPmos: -8.95199e+07 muA
** NormalTransistorNmos: 8.95191e+07 muA
** NormalTransistorNmos: 8.95181e+07 muA
** DiodeTransistorNmos: 1.78271e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.20801  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** inStageBiasComplementarySecondStage: 3.72501  V
** innerComplementarySecondStage: 2.98401  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.866001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.168001  V
** innerTransistorStack2Load1: 0.168001  V
** sourceTransconductance: 3.26801  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END