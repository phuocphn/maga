** Name: two_stage_single_output_op_amp_52_12

.MACRO two_stage_single_output_op_amp_52_12 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=70e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mMainBias3 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=92e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=14e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=93e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=30e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=6e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=70e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=44e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=44e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=268e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=93e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=120e-6
mMainBias15 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=72e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=492e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=307e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=307e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=553e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=267e-6
mMainBias21 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=76e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=600e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=492e-6
mMainBias24 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=345e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.2001e-12
.EOM two_stage_single_output_op_amp_52_12

** Expected Performance Values: 
** Gain: 172 dB
** Power consumption: 6.33901 mW
** Area: 14959 (mu_m)^2
** Transit frequency: 2.90101 MHz
** Transit frequency with error factor: 2.90089 MHz
** Slew rate: 3.62348 V/mu_s
** Phase margin: 63.0254°
** CMRR: 139 dB
** VoutMax: 4.25 V
** VoutMin: 1.29001 V
** VcmMax: 5.21001 V
** VcmMin: 0.810001 V


** Expected Currents: 
** NormalTransistorNmos: 2.03051e+07 muA
** NormalTransistorPmos: -1.16179e+08 muA
** NormalTransistorPmos: -8.98979e+07 muA
** NormalTransistorPmos: -2.55419e+07 muA
** NormalTransistorPmos: -6.66059e+07 muA
** NormalTransistorPmos: -1.04279e+08 muA
** NormalTransistorPmos: -6.66059e+07 muA
** NormalTransistorPmos: -1.04279e+08 muA
** DiodeTransistorNmos: 6.66051e+07 muA
** NormalTransistorNmos: 6.66051e+07 muA
** NormalTransistorNmos: 6.66051e+07 muA
** NormalTransistorNmos: 7.53451e+07 muA
** NormalTransistorNmos: 3.76731e+07 muA
** NormalTransistorNmos: 3.76731e+07 muA
** NormalTransistorNmos: 7.87323e+08 muA
** DiodeTransistorNmos: 7.87322e+08 muA
** NormalTransistorPmos: -7.87322e+08 muA
** NormalTransistorPmos: -7.87323e+08 muA
** DiodeTransistorNmos: 1.1618e+08 muA
** NormalTransistorNmos: 1.16179e+08 muA
** DiodeTransistorNmos: 8.98971e+07 muA
** DiodeTransistorNmos: 2.55411e+07 muA
** DiodeTransistorPmos: -2.03059e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.08301  V
** inputVoltageBiasXXnXX3: 0.587001  V
** out: 2.5  V
** outFirstStage: 4.15301  V
** outInputVoltageBiasXXnXX1: 1.70001  V
** outSourceVoltageBiasXXnXX1: 0.850001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.480001  V
** out1: 0.685001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.86901  V
** innerTransconductance: 4.71701  V
** inner: 0.850001  V


.END