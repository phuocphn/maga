** Name: two_stage_single_output_op_amp_26_1

.MACRO two_stage_single_output_op_amp_26_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=51e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=51e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=13e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=185e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=93e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=51e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=48e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=51e-6
mMainBias10 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=79e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=93e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=185e-6
mMainBias14 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mSecondStage1StageBias15 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=552e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.40001e-12
.EOM two_stage_single_output_op_amp_26_1

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 1.84101 mW
** Area: 3972 (mu_m)^2
** Transit frequency: 3.15601 MHz
** Transit frequency with error factor: 3.15109 MHz
** Slew rate: 5.9692 V/mu_s
** Phase margin: 60.1606°
** CMRR: 100 dB
** negPSRR: 95 dB
** posPSRR: 98 dB
** VoutMax: 4.84001 V
** VoutMin: 0.340001 V
** VcmMax: 3.18001 V
** VcmMin: 0.550001 V


** Expected Currents: 
** NormalTransistorNmos: 6.54561e+07 muA
** NormalTransistorPmos: -1.09599e+07 muA
** DiodeTransistorNmos: 1.61901e+07 muA
** NormalTransistorNmos: 1.61901e+07 muA
** NormalTransistorNmos: 1.61901e+07 muA
** DiodeTransistorNmos: 1.61901e+07 muA
** NormalTransistorPmos: -3.23829e+07 muA
** DiodeTransistorPmos: -3.23839e+07 muA
** NormalTransistorPmos: -1.61909e+07 muA
** NormalTransistorPmos: -1.61909e+07 muA
** NormalTransistorNmos: 2.39419e+08 muA
** NormalTransistorPmos: -2.39418e+08 muA
** DiodeTransistorNmos: 1.09591e+07 muA
** DiodeTransistorPmos: -6.54569e+07 muA
** NormalTransistorPmos: -6.54569e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.719001  V
** out: 2.5  V
** outFirstStage: 0.75  V
** outInputVoltageBiasXXpXX1: 3.47601  V
** outSourceVoltageBiasXXpXX1: 4.23801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.555001  V
** out1: 1.11001  V
** sourceTransconductance: 3.36401  V
** inner: 4.23801  V


.END