** Name: two_stage_single_output_op_amp_88_1

.MACRO two_stage_single_output_op_amp_88_1 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=136e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=10e-6 W=136e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=393e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=14e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=136e-6
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos4 L=10e-6 W=335e-6
mTelescopicFirstStageLoad8 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=136e-6
mMainBias9 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=189e-6
mTelescopicFirstStageLoad10 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=46e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=85e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=85e-6
mMainBias13 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=506e-6
mSecondStage1StageBias14 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=46e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=364e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.40001e-12
.EOM two_stage_single_output_op_amp_88_1

** Expected Performance Values: 
** Gain: 134 dB
** Power consumption: 3.20201 mW
** Area: 14418 (mu_m)^2
** Transit frequency: 3.64801 MHz
** Transit frequency with error factor: 3.64833 MHz
** Slew rate: 9.87511 V/mu_s
** Phase margin: 60.1606°
** CMRR: 136 dB
** VoutMax: 4.85001 V
** VoutMin: 0.300001 V
** VcmMax: 3.87001 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01997e+08 muA
** NormalTransistorPmos: -2.13806e+08 muA
** NormalTransistorPmos: -2.59039e+07 muA
** NormalTransistorPmos: -2.59039e+07 muA
** DiodeTransistorNmos: 2.59031e+07 muA
** DiodeTransistorNmos: 2.59031e+07 muA
** NormalTransistorNmos: 2.59031e+07 muA
** NormalTransistorNmos: 2.59031e+07 muA
** NormalTransistorPmos: -1.53805e+08 muA
** NormalTransistorPmos: -2.59049e+07 muA
** NormalTransistorPmos: -2.59049e+07 muA
** NormalTransistorNmos: 2.52694e+08 muA
** NormalTransistorPmos: -2.52693e+08 muA
** DiodeTransistorNmos: 2.13807e+08 muA
** DiodeTransistorPmos: -1.01996e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.565001  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outVoltageBiasXXpXX1: 2.27001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.47501  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 3.01101  V
** sourceGCC2: 3.01101  V


.END