** Name: two_stage_single_output_op_amp_21_3

.MACRO two_stage_single_output_op_amp_21_3 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=76e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=10e-6 W=57e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=19e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=76e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=437e-6
mSimpleFirstStageLoad7 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=10e-6 W=57e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=88e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=29e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=573e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=568e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=88e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_21_3

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 3.10101 mW
** Area: 7652 (mu_m)^2
** Transit frequency: 5.41801 MHz
** Transit frequency with error factor: 5.41405 MHz
** Slew rate: 6.69522 V/mu_s
** Phase margin: 69.9009°
** CMRR: 103 dB
** negPSRR: 99 dB
** posPSRR: 104 dB
** VoutMax: 3.96001 V
** VoutMin: 0.330001 V
** VcmMax: 3.20001 V
** VcmMin: 0.580001 V


** Expected Currents: 
** DiodeTransistorNmos: 1.52081e+07 muA
** DiodeTransistorNmos: 1.52071e+07 muA
** NormalTransistorNmos: 1.52081e+07 muA
** NormalTransistorNmos: 1.52071e+07 muA
** NormalTransistorPmos: -3.04169e+07 muA
** NormalTransistorPmos: -3.04159e+07 muA
** NormalTransistorPmos: -1.52089e+07 muA
** NormalTransistorPmos: -1.52089e+07 muA
** NormalTransistorNmos: 5.69794e+08 muA
** NormalTransistorPmos: -5.69793e+08 muA
** NormalTransistorPmos: -5.69794e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.46301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.735001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.558001  V
** innerStageBias: 4.26901  V
** innerTransistorStack2Load1: 0.557001  V
** out1: 1.14001  V
** sourceTransconductance: 3.26001  V
** innerStageBias: 4.26301  V


.END