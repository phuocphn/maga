** Name: two_stage_single_output_op_amp_177_5

.MACRO two_stage_single_output_op_amp_177_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=12e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=104e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=104e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=274e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=20e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=468e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=180e-6
mSimpleFirstStageLoad9 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=166e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=580e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=580e-6
mMainBias12 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=228e-6
mSecondStage1Transconductor13 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=55e-6
mSimpleFirstStageLoad14 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=166e-6
mMainBias15 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=52e-6
mSimpleFirstStageTransconductor16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=57e-6
mSimpleFirstStageStageBias17 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=41e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=104e-6
mSimpleFirstStageStageBias19 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=72e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=468e-6
mSimpleFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=104e-6
mSimpleFirstStageTransconductor23 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=57e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.90001e-12
.EOM two_stage_single_output_op_amp_177_5

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 6.33601 mW
** Area: 10932 (mu_m)^2
** Transit frequency: 3.41701 MHz
** Transit frequency with error factor: 3.41363 MHz
** Slew rate: 4.0674 V/mu_s
** Phase margin: 60.1606°
** CMRR: 122 dB
** VoutMax: 3.91001 V
** VoutMin: 0.700001 V
** VcmMax: 3.23001 V
** VcmMin: -0.129999 V


** Expected Currents: 
** NormalTransistorNmos: 2.47811e+07 muA
** NormalTransistorNmos: 1.08975e+08 muA
** DiodeTransistorPmos: -2.63988e+08 muA
** NormalTransistorPmos: -2.63987e+08 muA
** NormalTransistorPmos: -2.63988e+08 muA
** DiodeTransistorPmos: -2.63987e+08 muA
** NormalTransistorNmos: 2.76171e+08 muA
** NormalTransistorNmos: 2.76172e+08 muA
** NormalTransistorNmos: 2.76171e+08 muA
** NormalTransistorNmos: 2.76172e+08 muA
** NormalTransistorPmos: -2.43649e+07 muA
** NormalTransistorPmos: -2.43659e+07 muA
** NormalTransistorPmos: -1.21819e+07 muA
** NormalTransistorPmos: -1.21819e+07 muA
** NormalTransistorNmos: 5.71156e+08 muA
** NormalTransistorPmos: -5.71155e+08 muA
** DiodeTransistorPmos: -5.71156e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.47819e+07 muA
** NormalTransistorPmos: -2.47809e+07 muA
** DiodeTransistorPmos: -1.08974e+08 muA
** DiodeTransistorPmos: -1.08975e+08 muA


** Expected Voltages: 
** ibias: 1.15801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.40101  V
** out: 2.5  V
** outFirstStage: 1.10901  V
** outInputVoltageBiasXXpXX1: 3.34801  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.17401  V
** outSourceVoltageBiasXXpXX2: 4.17701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.74401  V
** innerSourceLoad1: 3.68601  V
** innerStageBias: 4.15901  V
** innerTransistorStack1Load1: 3.68401  V
** innerTransistorStack1Load2: 0.472001  V
** innerTransistorStack2Load2: 0.472001  V
** sourceTransconductance: 3.25301  V
** inner: 4.17501  V


.END