** Name: two_stage_single_output_op_amp_188_11

.MACRO two_stage_single_output_op_amp_188_11 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=74e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=9e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=105e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=20e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=102e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=201e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=42e-6
mSimpleFirstStageLoad9 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=74e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=20e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=509e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=105e-6
mSecondStage1StageBias13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=528e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=89e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=42e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=526e-6
mMainBias17 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=250e-6
mSimpleFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=587e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=586e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=269e-6
mSimpleFirstStageLoad21 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=587e-6
mMainBias22 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=113e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_188_11

** Expected Performance Values: 
** Gain: 110 dB
** Power consumption: 14.3311 mW
** Area: 14943 (mu_m)^2
** Transit frequency: 6.03701 MHz
** Transit frequency with error factor: 5.89218 MHz
** Slew rate: 5.6899 V/mu_s
** Phase margin: 66.4632°
** CMRR: 97 dB
** VoutMax: 4.32001 V
** VoutMin: 0.710001 V
** VcmMax: 4.82001 V
** VcmMin: 1.46001 V


** Expected Currents: 
** NormalTransistorNmos: 5.17823e+08 muA
** NormalTransistorNmos: 2.45246e+08 muA
** NormalTransistorPmos: -1.40282e+08 muA
** NormalTransistorNmos: 7.11676e+08 muA
** NormalTransistorNmos: 7.11677e+08 muA
** DiodeTransistorNmos: 7.11676e+08 muA
** NormalTransistorPmos: -7.25008e+08 muA
** NormalTransistorPmos: -7.25008e+08 muA
** NormalTransistorNmos: 2.66651e+07 muA
** DiodeTransistorNmos: 2.66641e+07 muA
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 5.02823e+08 muA
** NormalTransistorNmos: 5.02822e+08 muA
** NormalTransistorPmos: -5.02822e+08 muA
** NormalTransistorPmos: -5.02823e+08 muA
** DiodeTransistorNmos: 1.40283e+08 muA
** NormalTransistorNmos: 1.40282e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.17822e+08 muA
** DiodeTransistorPmos: -2.45245e+08 muA


** Expected Voltages: 
** ibias: 1.125  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.21601  V
** outInputVoltageBiasXXnXX1: 1.31001  V
** outSourceVoltageBiasXXnXX1: 0.655001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 3.84901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.570001  V
** innerTransconductance: 4.70601  V
** inner: 0.653001  V


.END