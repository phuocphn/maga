** Name: two_stage_single_output_op_amp_78_11

.MACRO two_stage_single_output_op_amp_78_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=7e-6 W=24e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=26e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=8e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=194e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=90e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=5e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=386e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=26e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=18e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=18e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=90e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=546e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=194e-6
mSecondStage1StageBias15 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=569e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=24e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=99e-6
mFoldedCascodeFirstStageLoad19 FirstStageYinnerOutputLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=108e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=103e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=103e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=546e-6
mSecondStage1Transconductor23 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=348e-6
mFoldedCascodeFirstStageLoad24 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=108e-6
mMainBias25 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=150e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_78_11

** Expected Performance Values: 
** Gain: 177 dB
** Power consumption: 3.77301 mW
** Area: 14985 (mu_m)^2
** Transit frequency: 4.00601 MHz
** Transit frequency with error factor: 4.00614 MHz
** Slew rate: 3.77575 V/mu_s
** Phase margin: 64.1713°
** CMRR: 144 dB
** VoutMax: 4.26001 V
** VoutMin: 0.710001 V
** VcmMax: 5.14001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 1.69211e+07 muA
** NormalTransistorNmos: 9.71171e+07 muA
** NormalTransistorPmos: -3.73239e+07 muA
** NormalTransistorPmos: -1.71429e+07 muA
** NormalTransistorPmos: -2.57129e+07 muA
** NormalTransistorPmos: -1.71469e+07 muA
** NormalTransistorPmos: -2.57189e+07 muA
** DiodeTransistorNmos: 1.71441e+07 muA
** DiodeTransistorNmos: 1.71451e+07 muA
** NormalTransistorNmos: 1.71461e+07 muA
** NormalTransistorNmos: 1.71451e+07 muA
** NormalTransistorNmos: 1.71421e+07 muA
** DiodeTransistorNmos: 1.71421e+07 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 5.41867e+08 muA
** NormalTransistorNmos: 5.41866e+08 muA
** NormalTransistorPmos: -5.41866e+08 muA
** NormalTransistorPmos: -5.41867e+08 muA
** DiodeTransistorNmos: 3.73231e+07 muA
** NormalTransistorNmos: 3.73221e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.69219e+07 muA
** DiodeTransistorPmos: -9.71179e+07 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.20001  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.17101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.28501  V
** innerTransistorStack1Load2: 0.638001  V
** innerTransistorStack2Load2: 0.636001  V
** sourceGCC1: 4.41301  V
** sourceGCC2: 4.41301  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.579001  V
** innerTransconductance: 4.75901  V
** inner: 0.554001  V


.END