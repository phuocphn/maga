** Name: two_stage_single_output_op_amp_19_1

.MACRO two_stage_single_output_op_amp_19_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=30e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=11e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=36e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=10e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=30e-6
mMainBias7 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=227e-6
mSimpleFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=23e-6
mSimpleFirstStageTransconductor10 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=59e-6
mSimpleFirstStageStageBias11 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=58e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=8e-6 W=90e-6
mMainBias13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=29e-6
mSecondStage1StageBias14 out ibias sourcePmos sourcePmos pmos4 L=4e-6 W=512e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=59e-6
mMainBias16 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=25e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_19_1

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 1.01001 mW
** Area: 5279 (mu_m)^2
** Transit frequency: 3.77201 MHz
** Transit frequency with error factor: 3.7694 MHz
** Slew rate: 3.61195 V/mu_s
** Phase margin: 65.3172°
** CMRR: 106 dB
** negPSRR: 108 dB
** posPSRR: 215 dB
** VoutMax: 4.75 V
** VoutMin: 0.150001 V
** VcmMax: 3.19001 V
** VcmMin: 0.150001 V


** Expected Currents: 
** NormalTransistorNmos: 6.41901e+06 muA
** NormalTransistorPmos: -7.04999e+06 muA
** NormalTransistorPmos: -8.11199e+06 muA
** DiodeTransistorNmos: 8.16301e+06 muA
** NormalTransistorNmos: 8.16301e+06 muA
** NormalTransistorNmos: 8.16301e+06 muA
** NormalTransistorPmos: -1.63269e+07 muA
** NormalTransistorPmos: -1.63279e+07 muA
** NormalTransistorPmos: -8.16399e+06 muA
** NormalTransistorPmos: -8.16399e+06 muA
** NormalTransistorNmos: 1.4414e+08 muA
** NormalTransistorPmos: -1.44139e+08 muA
** DiodeTransistorNmos: 7.04901e+06 muA
** DiodeTransistorNmos: 8.11101e+06 muA
** DiodeTransistorPmos: -6.41999e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.713001  V
** inputVoltageBiasXXpXX1: 3.89801  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.679001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerStageBias: 4.74601  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.21601  V


.END