** Name: two_stage_single_output_op_amp_34_9

.MACRO two_stage_single_output_op_amp_34_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=34e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=319e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=333e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=555e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
mMainBias7 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=25e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=319e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=34e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mMainBias13 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mSecondStage1StageBias14 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=333e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=25e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=555e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad18 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=497e-6
mMainBias19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=56e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.90001e-12
.EOM two_stage_single_output_op_amp_34_9

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 6.22901 mW
** Area: 7739 (mu_m)^2
** Transit frequency: 9.32101 MHz
** Transit frequency with error factor: 9.29408 MHz
** Slew rate: 22.6166 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** negPSRR: 134 dB
** posPSRR: 90 dB
** VoutMax: 4.75 V
** VoutMin: 0.840001 V
** VcmMax: 4.44001 V
** VcmMin: 1.90001 V


** Expected Currents: 
** NormalTransistorNmos: 3.42231e+07 muA
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -4.21529e+07 muA
** DiodeTransistorPmos: -1.99947e+08 muA
** NormalTransistorPmos: -1.99947e+08 muA
** NormalTransistorPmos: -1.99947e+08 muA
** NormalTransistorNmos: 3.99894e+08 muA
** DiodeTransistorNmos: 3.99893e+08 muA
** NormalTransistorNmos: 1.99948e+08 muA
** NormalTransistorNmos: 1.99948e+08 muA
** NormalTransistorNmos: 6.58087e+08 muA
** DiodeTransistorNmos: 6.58086e+08 muA
** NormalTransistorPmos: -6.58086e+08 muA
** DiodeTransistorNmos: 4.21521e+07 muA
** NormalTransistorNmos: 4.21521e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.42239e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 1.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.23101  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.18901  V
** outInputVoltageBiasXXnXX1: 1.15401  V
** outSourceVoltageBiasXXnXX1: 0.577001  V
** outSourceVoltageBiasXXnXX2: 0.622001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.40001  V
** out1: 4.18901  V
** sourceTransconductance: 1.34501  V
** inner: 0.577001  V
** inner: 0.619001  V


.END