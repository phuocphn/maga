** Name: two_stage_single_output_op_amp_188_9

.MACRO two_stage_single_output_op_amp_188_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=10e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=6e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=7e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=60e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=271e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=47e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=10e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=60e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=271e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=8e-6 W=19e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=47e-6
mSimpleFirstStageLoad15 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=224e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=527e-6
mSimpleFirstStageLoad17 outFirstStage ibias sourcePmos sourcePmos pmos4 L=3e-6 W=224e-6
mMainBias18 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=18e-6
mMainBias19 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=136e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.1001e-12
.EOM two_stage_single_output_op_amp_188_9

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 14.9931 mW
** Area: 5888 (mu_m)^2
** Transit frequency: 6.26101 MHz
** Transit frequency with error factor: 6.2525 MHz
** Slew rate: 5.90123 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 1.76001 V
** VcmMax: 5.11001 V
** VcmMin: 1.33001 V


** Expected Currents: 
** NormalTransistorPmos: -9.06799e+06 muA
** NormalTransistorPmos: -6.79609e+07 muA
** NormalTransistorNmos: 6.83541e+07 muA
** NormalTransistorNmos: 6.83551e+07 muA
** DiodeTransistorNmos: 6.83541e+07 muA
** NormalTransistorPmos: -1.13113e+08 muA
** NormalTransistorPmos: -1.13113e+08 muA
** NormalTransistorNmos: 8.95171e+07 muA
** DiodeTransistorNmos: 8.95161e+07 muA
** NormalTransistorNmos: 4.47591e+07 muA
** NormalTransistorNmos: 4.47591e+07 muA
** NormalTransistorNmos: 2.67543e+09 muA
** DiodeTransistorNmos: 2.67543e+09 muA
** NormalTransistorPmos: -2.67542e+09 muA
** DiodeTransistorNmos: 9.06701e+06 muA
** NormalTransistorNmos: 9.06601e+06 muA
** DiodeTransistorNmos: 6.79601e+07 muA
** NormalTransistorNmos: 6.79591e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.14501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.18501  V
** outInputVoltageBiasXXnXX2: 2.17001  V
** outSourceVoltageBiasXXnXX1: 0.593001  V
** outSourceVoltageBiasXXnXX2: 1.08501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** out1: 2.14601  V
** sourceTransconductance: 1.94501  V
** inner: 0.591001  V
** inner: 1.08501  V


.END