** Name: two_stage_single_output_op_amp_133_1

.MACRO two_stage_single_output_op_amp_133_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=46e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=46e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mSimpleFirstStageLoad5 FirstStageYinnerOutputLoad1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=94e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=458e-6
mSimpleFirstStageLoad7 outFirstStage outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=94e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=56e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=46e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=310e-6
mSecondStage1StageBias11 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=46e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=56e-6
mMainBias14 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.7001e-12
.EOM two_stage_single_output_op_amp_133_1

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 3.98601 mW
** Area: 3725 (mu_m)^2
** Transit frequency: 4.18601 MHz
** Transit frequency with error factor: 4.1664 MHz
** Slew rate: 8.34258 V/mu_s
** Phase margin: 60.1606°
** CMRR: 80 dB
** VoutMax: 4.84001 V
** VoutMin: 0.150001 V
** VcmMax: 3.89001 V
** VcmMin: -0.269999 V


** Expected Currents: 
** NormalTransistorPmos: -2.41489e+07 muA
** DiodeTransistorPmos: -1.55684e+08 muA
** DiodeTransistorPmos: -1.55684e+08 muA
** NormalTransistorPmos: -1.55684e+08 muA
** NormalTransistorPmos: -1.55684e+08 muA
** NormalTransistorNmos: 2.30918e+08 muA
** NormalTransistorNmos: 2.30918e+08 muA
** NormalTransistorPmos: -1.50466e+08 muA
** NormalTransistorPmos: -7.52329e+07 muA
** NormalTransistorPmos: -7.52329e+07 muA
** NormalTransistorNmos: 2.91288e+08 muA
** NormalTransistorPmos: -2.91287e+08 muA
** DiodeTransistorNmos: 2.41481e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX1: 0.699001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerSourceLoad1: 3.68601  V
** innerTransistorStack2Load1: 3.68601  V
** sourceTransconductance: 3.45001  V


.END