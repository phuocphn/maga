** Name: two_stage_single_output_op_amp_162_3

.MACRO two_stage_single_output_op_amp_162_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=40e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=47e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=12e-6
mMainBias5 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=3e-6 W=4e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=168e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=183e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=183e-6
mSimpleFirstStageLoad10 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=173e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=94e-6
mSimpleFirstStageLoad12 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=173e-6
mMainBias13 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mMainBias14 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=51e-6
mSimpleFirstStageTransconductor15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=44e-6
mSimpleFirstStageLoad16 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSimpleFirstStageStageBias17 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=168e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=288e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=12e-6
mSecondStage1StageBias20 out outInputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=246e-6
mSimpleFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=10e-6 W=25e-6
mSimpleFirstStageTransconductor22 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=44e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.20001e-12
.EOM two_stage_single_output_op_amp_162_3

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 4.36101 mW
** Area: 12145 (mu_m)^2
** Transit frequency: 3.55601 MHz
** Transit frequency with error factor: 3.55477 MHz
** Slew rate: 5.04202 V/mu_s
** Phase margin: 60.1606°
** CMRR: 94 dB
** VoutMax: 3.04001 V
** VoutMin: 0.310001 V
** VcmMax: 3.18001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 1.90501e+06 muA
** NormalTransistorNmos: 1.09011e+07 muA
** NormalTransistorPmos: -2.53829e+07 muA
** NormalTransistorPmos: -2.53829e+07 muA
** DiodeTransistorPmos: -2.53829e+07 muA
** NormalTransistorNmos: 3.87271e+07 muA
** NormalTransistorNmos: 3.87281e+07 muA
** NormalTransistorNmos: 3.87271e+07 muA
** NormalTransistorNmos: 3.87281e+07 muA
** NormalTransistorPmos: -2.66909e+07 muA
** DiodeTransistorPmos: -2.66919e+07 muA
** NormalTransistorPmos: -1.33449e+07 muA
** NormalTransistorPmos: -1.33449e+07 muA
** NormalTransistorNmos: 7.71832e+08 muA
** NormalTransistorPmos: -7.71831e+08 muA
** NormalTransistorPmos: -7.71832e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.90599e+06 muA
** NormalTransistorPmos: -1.90699e+06 muA
** DiodeTransistorPmos: -1.09019e+07 muA
** DiodeTransistorPmos: -1.09029e+07 muA


** Expected Voltages: 
** ibias: 1.12301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.718001  V
** outInputVoltageBiasXXpXX1: 3.40801  V
** outInputVoltageBiasXXpXX2: 2.51901  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.20401  V
** outSourceVoltageBiasXXpXX2: 3.76201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.68601  V
** innerTransistorStack1Load2: 0.563001  V
** innerTransistorStack2Load2: 0.563001  V
** out1: 2.37201  V
** sourceTransconductance: 3.28901  V
** innerStageBias: 3.80601  V
** inner: 4.20201  V


.END