** Name: two_stage_single_output_op_amp_72_1

.MACRO two_stage_single_output_op_amp_72_1 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=97e-6
mMainBias2 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=13e-6
mFoldedCascodeFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=83e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=14e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
mFoldedCascodeFirstStageTransconductor6 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=55e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=55e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=83e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=13e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=587e-6
mFoldedCascodeFirstStageLoad11 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=97e-6
mMainBias12 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=37e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=112e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=5e-6 W=588e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mSecondStage1StageBias17 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=564e-6
mFoldedCascodeFirstStageLoad18 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=5e-6 W=588e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.5e-12
.EOM two_stage_single_output_op_amp_72_1

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 7.00701 mW
** Area: 10706 (mu_m)^2
** Transit frequency: 3.64901 MHz
** Transit frequency with error factor: 3.64819 MHz
** Slew rate: 3.50356 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** VoutMax: 4.67001 V
** VoutMin: 0.150001 V
** VcmMax: 5.07001 V
** VcmMin: 1.48001 V


** Expected Currents: 
** NormalTransistorNmos: 2.84281e+07 muA
** NormalTransistorNmos: 8.65851e+07 muA
** NormalTransistorPmos: -4.77609e+07 muA
** NormalTransistorPmos: -7.92329e+07 muA
** NormalTransistorPmos: -4.77609e+07 muA
** NormalTransistorPmos: -7.92329e+07 muA
** DiodeTransistorNmos: 4.77601e+07 muA
** NormalTransistorNmos: 4.77601e+07 muA
** NormalTransistorNmos: 6.29421e+07 muA
** DiodeTransistorNmos: 6.29431e+07 muA
** NormalTransistorNmos: 3.14711e+07 muA
** NormalTransistorNmos: 3.14711e+07 muA
** NormalTransistorNmos: 1.11802e+09 muA
** NormalTransistorPmos: -1.11801e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.84289e+07 muA
** DiodeTransistorPmos: -8.65859e+07 muA


** Expected Voltages: 
** ibias: 1.27401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXnXX1: 0.638001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.10201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.557001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.89301  V
** inner: 0.635001  V


.END