** Name: two_stage_single_output_op_amp_11_9

.MACRO two_stage_single_output_op_amp_11_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=11e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=269e-6
mSimpleFirstStageLoad4 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=8e-6 W=158e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=33e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=14e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=12e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=14e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mSecondStage1StageBias10 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=269e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=12e-6
mMainBias12 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=33e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=205e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=8e-6 W=158e-6
mMainBias16 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=30e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_11_9

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 2.90401 mW
** Area: 5164 (mu_m)^2
** Transit frequency: 2.92001 MHz
** Transit frequency with error factor: 2.91584 MHz
** Slew rate: 6.03322 V/mu_s
** Phase margin: 63.5984°
** CMRR: 101 dB
** negPSRR: 92 dB
** posPSRR: 87 dB
** VoutMax: 4.25 V
** VoutMin: 0.700001 V
** VcmMax: 3.65001 V
** VcmMin: 1.04001 V


** Expected Currents: 
** NormalTransistorNmos: 9.96501e+06 muA
** NormalTransistorPmos: -2.09519e+07 muA
** DiodeTransistorPmos: -1.37349e+07 muA
** DiodeTransistorPmos: -1.37359e+07 muA
** NormalTransistorPmos: -1.37349e+07 muA
** NormalTransistorPmos: -1.37359e+07 muA
** NormalTransistorNmos: 2.74681e+07 muA
** NormalTransistorNmos: 1.37341e+07 muA
** NormalTransistorNmos: 1.37341e+07 muA
** NormalTransistorNmos: 5.12346e+08 muA
** DiodeTransistorNmos: 5.12346e+08 muA
** NormalTransistorPmos: -5.12345e+08 muA
** DiodeTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.96599e+06 muA


** Expected Voltages: 
** ibias: 0.711001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX0: 3.80801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.24101  V
** innerSourceLoad1: 4.00301  V
** innerTransistorStack2Load1: 4.00201  V
** sourceTransconductance: 1.76501  V
** inner: 0.555001  V


.END