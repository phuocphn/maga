** Name: two_stage_single_output_op_amp_53_11

.MACRO two_stage_single_output_op_amp_53_11 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=145e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=5e-6 W=338e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mMainBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=23e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=93e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=145e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=20e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=20e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=136e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=463e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=416e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=338e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=62e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=30e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=150e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=555e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=555e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=521e-6
mMainBias20 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=324e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=600e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=150e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.5e-12
.EOM two_stage_single_output_op_amp_53_11

** Expected Performance Values: 
** Gain: 156 dB
** Power consumption: 6.44501 mW
** Area: 14960 (mu_m)^2
** Transit frequency: 2.92001 MHz
** Transit frequency with error factor: 2.91951 MHz
** Slew rate: 9.20579 V/mu_s
** Phase margin: 61.3065°
** CMRR: 128 dB
** VoutMax: 4.25 V
** VoutMin: 0.5 V
** VcmMax: 5.25 V
** VcmMin: 1.24001 V


** Expected Currents: 
** NormalTransistorNmos: 7.76161e+07 muA
** NormalTransistorNmos: 3.75561e+07 muA
** NormalTransistorPmos: -1.32329e+08 muA
** NormalTransistorPmos: -1.43681e+08 muA
** NormalTransistorPmos: -2.2842e+08 muA
** NormalTransistorPmos: -1.43681e+08 muA
** NormalTransistorPmos: -2.2842e+08 muA
** DiodeTransistorNmos: 1.43682e+08 muA
** DiodeTransistorNmos: 1.43681e+08 muA
** NormalTransistorNmos: 1.43682e+08 muA
** NormalTransistorNmos: 1.43681e+08 muA
** NormalTransistorNmos: 1.69476e+08 muA
** NormalTransistorNmos: 8.47381e+07 muA
** NormalTransistorNmos: 8.47381e+07 muA
** NormalTransistorNmos: 5.74731e+08 muA
** NormalTransistorNmos: 5.7473e+08 muA
** NormalTransistorPmos: -5.7473e+08 muA
** NormalTransistorPmos: -5.74731e+08 muA
** DiodeTransistorNmos: 1.3233e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.76169e+07 muA
** DiodeTransistorPmos: -3.75569e+07 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.10201  V
** out: 2.5  V
** outFirstStage: 4.08501  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.28501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.646001  V
** innerTransistorStack2Load2: 0.645001  V
** out1: 1.20901  V
** sourceGCC1: 4.64901  V
** sourceGCC2: 4.64901  V
** sourceTransconductance: 1.50101  V
** innerStageBias: 0.442001  V
** innerTransconductance: 4.64901  V


.END