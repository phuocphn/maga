** Name: two_stage_single_output_op_amp_130_4

.MACRO two_stage_single_output_op_amp_130_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=9e-6 W=89e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=18e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=113e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=113e-6
mSimpleFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=55e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=522e-6
mMainBias10 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=120e-6
mSecondStage1Transconductor11 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=347e-6
mSimpleFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=55e-6
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=341e-6
mSimpleFirstStageLoad14 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=9e-6 W=89e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=228e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=594e-6
mMainBias17 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=229e-6
mMainBias18 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=74e-6
mSecondStage1StageBias19 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=599e-6
mSimpleFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=5e-6 W=49e-6
mSimpleFirstStageTransconductor21 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=341e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.6001e-12
.EOM two_stage_single_output_op_amp_130_4

** Expected Performance Values: 
** Gain: 148 dB
** Power consumption: 5.12601 mW
** Area: 14977 (mu_m)^2
** Transit frequency: 3.57501 MHz
** Transit frequency with error factor: 3.57169 MHz
** Slew rate: 6.52215 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.52001 V
** VoutMin: 0.300001 V
** VcmMax: 3.84001 V
** VcmMin: -0.0699999 V


** Expected Currents: 
** NormalTransistorNmos: 1.72607e+08 muA
** NormalTransistorPmos: -1.29015e+08 muA
** NormalTransistorPmos: -4.13819e+07 muA
** NormalTransistorPmos: -9.95039e+07 muA
** NormalTransistorPmos: -9.95029e+07 muA
** DiodeTransistorPmos: -9.95039e+07 muA
** NormalTransistorNmos: 1.63731e+08 muA
** NormalTransistorNmos: 1.6373e+08 muA
** NormalTransistorNmos: 1.6373e+08 muA
** NormalTransistorNmos: 1.6373e+08 muA
** NormalTransistorPmos: -1.28452e+08 muA
** NormalTransistorPmos: -6.42269e+07 muA
** NormalTransistorPmos: -6.42269e+07 muA
** NormalTransistorNmos: 3.34654e+08 muA
** NormalTransistorNmos: 3.34653e+08 muA
** NormalTransistorPmos: -3.34653e+08 muA
** NormalTransistorPmos: -3.34654e+08 muA
** DiodeTransistorNmos: 1.29016e+08 muA
** DiodeTransistorNmos: 4.13811e+07 muA
** DiodeTransistorPmos: -1.72606e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.907001  V
** inputVoltageBiasXXnXX2: 0.631001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.236001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.236001  V
** out1: 2.37201  V
** sourceTransconductance: 3.35301  V
** innerStageBias: 4.42601  V
** innerTransconductance: 0.351001  V


.END