** Name: two_stage_single_output_op_amp_23_4

.MACRO two_stage_single_output_op_amp_23_4 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=49e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=13e-6
mMainBias3 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=63e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=143e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=143e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=280e-6
mSecondStage1Transconductor8 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=464e-6
mSimpleFirstStageLoad9 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=63e-6
mSimpleFirstStageTransconductor10 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=498e-6
mSimpleFirstStageStageBias11 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=120e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=79e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=529e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=344e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=498e-6
mMainBias16 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=271e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.20001e-12
.EOM two_stage_single_output_op_amp_23_4

** Expected Performance Values: 
** Gain: 148 dB
** Power consumption: 4.76401 mW
** Area: 11474 (mu_m)^2
** Transit frequency: 11.4931 MHz
** Transit frequency with error factor: 11.4833 MHz
** Slew rate: 14.6246 V/mu_s
** Phase margin: 60.1606°
** CMRR: 101 dB
** negPSRR: 105 dB
** posPSRR: 124 dB
** VoutMax: 3.91001 V
** VoutMin: 0.320001 V
** VcmMax: 3.14001 V
** VcmMin: -0.349999 V


** Expected Currents: 
** NormalTransistorPmos: -2.7476e+08 muA
** NormalTransistorNmos: 6.08321e+07 muA
** NormalTransistorNmos: 6.08311e+07 muA
** NormalTransistorNmos: 6.08321e+07 muA
** NormalTransistorNmos: 6.08311e+07 muA
** NormalTransistorPmos: -1.21665e+08 muA
** NormalTransistorPmos: -1.21664e+08 muA
** NormalTransistorPmos: -6.08329e+07 muA
** NormalTransistorPmos: -6.08329e+07 muA
** NormalTransistorNmos: 5.36342e+08 muA
** NormalTransistorNmos: 5.36341e+08 muA
** NormalTransistorPmos: -5.36341e+08 muA
** NormalTransistorPmos: -5.3634e+08 muA
** DiodeTransistorNmos: 2.74761e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.42701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.768001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.617001  V
** innerStageBias: 4.28401  V
** innerTransistorStack1Load1: 0.212001  V
** innerTransistorStack2Load1: 0.212001  V
** sourceTransconductance: 3.26601  V
** innerStageBias: 4.28501  V
** innerTransconductance: 0.197001  V


.END