** Name: two_stage_single_output_op_amp_71_4

.MACRO two_stage_single_output_op_amp_71_4 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=16e-6
mSecondStage1StageBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=34e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=95e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=21e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=15e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=29e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=12e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=234e-6
mSecondStage1Transconductor11 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=170e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=16e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=320e-6
mMainBias17 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=235e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=99e-6
mSecondStage1StageBias19 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=596e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=39e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_71_4

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 3.63601 mW
** Area: 5313 (mu_m)^2
** Transit frequency: 3.48501 MHz
** Transit frequency with error factor: 3.48076 MHz
** Slew rate: 3.52408 V/mu_s
** Phase margin: 62.4525°
** CMRR: 102 dB
** VoutMax: 4.03001 V
** VoutMin: 0.700001 V
** VcmMax: 5.17001 V
** VcmMin: 1.44001 V


** Expected Currents: 
** NormalTransistorPmos: -2.34717e+08 muA
** NormalTransistorPmos: -1.00372e+08 muA
** NormalTransistorPmos: -1.59029e+07 muA
** NormalTransistorPmos: -2.38529e+07 muA
** NormalTransistorPmos: -1.59049e+07 muA
** NormalTransistorPmos: -2.38569e+07 muA
** DiodeTransistorNmos: 1.59041e+07 muA
** NormalTransistorNmos: 1.59041e+07 muA
** NormalTransistorNmos: 1.59011e+07 muA
** NormalTransistorNmos: 1.59001e+07 muA
** NormalTransistorNmos: 7.95101e+06 muA
** NormalTransistorNmos: 7.95101e+06 muA
** NormalTransistorNmos: 3.24442e+08 muA
** NormalTransistorNmos: 3.24441e+08 muA
** NormalTransistorPmos: -3.24441e+08 muA
** NormalTransistorPmos: -3.2444e+08 muA
** DiodeTransistorNmos: 2.34718e+08 muA
** DiodeTransistorNmos: 1.00373e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.10801  V
** inputVoltageBiasXXnXX2: 0.563001  V
** out: 2.5  V
** outFirstStage: 0.742001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.729001  V
** innerStageBias: 0.396001  V
** sourceGCC1: 4.18601  V
** sourceGCC2: 4.18601  V
** sourceTransconductance: 1.93401  V
** innerStageBias: 4.20901  V
** innerTransconductance: 0.337001  V


.END