** Name: two_stage_single_output_op_amp_31_12

.MACRO two_stage_single_output_op_amp_31_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=14e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=312e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=3e-6 W=398e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=64e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=175e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=61e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=181e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=312e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=61e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=367e-6
mSimpleFirstStageLoad16 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=3e-6 W=398e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=511e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=93e-6
mMainBias20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=208e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.4001e-12
.EOM two_stage_single_output_op_amp_31_12

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 9.26101 mW
** Area: 11447 (mu_m)^2
** Transit frequency: 9.90601 MHz
** Transit frequency with error factor: 9.90074 MHz
** Slew rate: 9.336 V/mu_s
** Phase margin: 60.1606°
** CMRR: 108 dB
** negPSRR: 107 dB
** posPSRR: 100 dB
** VoutMax: 4.25 V
** VoutMin: 1.53001 V
** VcmMax: 4.5 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 1.92961e+07 muA
** NormalTransistorNmos: 2.43681e+08 muA
** NormalTransistorPmos: -6.17679e+07 muA
** NormalTransistorPmos: -5.80929e+07 muA
** NormalTransistorPmos: -5.80929e+07 muA
** DiodeTransistorPmos: -5.80929e+07 muA
** NormalTransistorNmos: 1.16184e+08 muA
** NormalTransistorNmos: 1.16183e+08 muA
** NormalTransistorNmos: 5.80921e+07 muA
** NormalTransistorNmos: 5.80921e+07 muA
** NormalTransistorNmos: 1.40127e+09 muA
** DiodeTransistorNmos: 1.40127e+09 muA
** NormalTransistorPmos: -1.40126e+09 muA
** NormalTransistorPmos: -1.40126e+09 muA
** DiodeTransistorNmos: 6.17671e+07 muA
** NormalTransistorNmos: 6.17671e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.92969e+07 muA
** DiodeTransistorPmos: -2.4368e+08 muA


** Expected Voltages: 
** ibias: 1.22801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.14701  V
** out: 2.5  V
** outFirstStage: 4.04601  V
** outInputVoltageBiasXXnXX1: 1.93401  V
** outSourceVoltageBiasXXnXX1: 0.967001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.672001  V
** innerTransistorStack2Load1: 4.28001  V
** out1: 3.52901  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.61001  V
** inner: 0.967001  V


.END