** Name: two_stage_single_output_op_amp_46_5

.MACRO two_stage_single_output_op_amp_46_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=5e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=286e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=7e-6 W=61e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=5e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=251e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=282e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=7e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=106e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=7e-6
mMainBias13 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=17e-6
mMainBias14 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=46e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=286e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=104e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=104e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=167e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
mSecondStage1StageBias20 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=251e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=61e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_46_5

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 3.34601 mW
** Area: 10909 (mu_m)^2
** Transit frequency: 4.03201 MHz
** Transit frequency with error factor: 4.03212 MHz
** Slew rate: 3.84794 V/mu_s
** Phase margin: 61.3065°
** CMRR: 136 dB
** VoutMax: 3.01001 V
** VoutMin: 0.620001 V
** VcmMax: 4.13001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.12421e+07 muA
** NormalTransistorNmos: 3.00841e+07 muA
** NormalTransistorNmos: 1.73671e+07 muA
** NormalTransistorNmos: 2.61601e+07 muA
** NormalTransistorNmos: 1.73671e+07 muA
** NormalTransistorNmos: 2.61601e+07 muA
** DiodeTransistorPmos: -1.73679e+07 muA
** DiodeTransistorPmos: -1.73689e+07 muA
** NormalTransistorPmos: -1.73679e+07 muA
** NormalTransistorPmos: -1.73689e+07 muA
** NormalTransistorPmos: -1.75889e+07 muA
** NormalTransistorPmos: -8.79399e+06 muA
** NormalTransistorPmos: -8.79399e+06 muA
** NormalTransistorNmos: 5.65507e+08 muA
** NormalTransistorPmos: -5.65506e+08 muA
** DiodeTransistorPmos: -5.65507e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.12429e+07 muA
** NormalTransistorPmos: -1.12439e+07 muA
** DiodeTransistorPmos: -3.00849e+07 muA


** Expected Voltages: 
** ibias: 1.22801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 1.02301  V
** outInputVoltageBiasXXpXX1: 2.44601  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 3.72301  V
** outVoltageBiasXXpXX2: 4.28201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.28101  V
** innerTransistorStack2Load2: 4.27901  V
** out1: 3.38201  V
** sourceGCC1: 0.525001  V
** sourceGCC2: 0.525001  V
** sourceTransconductance: 3.21801  V
** inner: 3.71601  V


.END