** Name: two_stage_single_output_op_amp_118_8

.MACRO two_stage_single_output_op_amp_118_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=4e-6 W=8e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=11e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=23e-6
mTelescopicFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=41e-6
mMainBias5 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=73e-6
mMainBias7 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=23e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=8e-6
mTelescopicFirstStageLoad9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=75e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=75e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=75e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=152e-6
mTelescopicFirstStageLoad15 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=75e-6
mMainBias16 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=41e-6
mTelescopicFirstStageStageBias18 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=41e-6
mTelescopicFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=73e-6
mMainBias20 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=48e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=538e-6
mTelescopicFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=203e-6
mMainBias23 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=117e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.4001e-12
.EOM two_stage_single_output_op_amp_118_8

** Expected Performance Values: 
** Gain: 154 dB
** Power consumption: 2.03001 mW
** Area: 10541 (mu_m)^2
** Transit frequency: 2.98901 MHz
** Transit frequency with error factor: 2.98943 MHz
** Slew rate: 3.63573 V/mu_s
** Phase margin: 60.1606°
** CMRR: 147 dB
** VoutMax: 4.83001 V
** VoutMin: 0.850001 V
** VcmMax: 4.16001 V
** VcmMin: 1.51001 V


** Expected Currents: 
** NormalTransistorNmos: 5.77101e+06 muA
** NormalTransistorNmos: 1.96611e+07 muA
** NormalTransistorPmos: -2.94059e+07 muA
** NormalTransistorPmos: -1.18549e+07 muA
** NormalTransistorNmos: 2.04071e+07 muA
** NormalTransistorNmos: 2.04071e+07 muA
** DiodeTransistorPmos: -2.04079e+07 muA
** NormalTransistorPmos: -2.04079e+07 muA
** NormalTransistorPmos: -2.04079e+07 muA
** NormalTransistorNmos: 5.26671e+07 muA
** DiodeTransistorNmos: 5.26661e+07 muA
** NormalTransistorNmos: 2.04071e+07 muA
** NormalTransistorNmos: 2.04071e+07 muA
** NormalTransistorNmos: 2.88581e+08 muA
** NormalTransistorNmos: 2.8858e+08 muA
** NormalTransistorPmos: -2.8858e+08 muA
** DiodeTransistorNmos: 2.94051e+07 muA
** NormalTransistorNmos: 2.94041e+07 muA
** DiodeTransistorNmos: 1.18541e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -5.77199e+06 muA
** DiodeTransistorPmos: -1.96619e+07 muA


** Expected Voltages: 
** ibias: 1.20201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 2.65001  V
** out: 2.5  V
** outFirstStage: 4.26201  V
** outInputVoltageBiasXXnXX1: 1.36001  V
** outSourceVoltageBiasXXnXX1: 0.680001  V
** outSourceVoltageBiasXXnXX3: 0.555001  V
** outVoltageBiasXXpXX0: 4.08201  V
** outVoltageBiasXXpXX1: 3.69801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 4.41201  V
** out1: 4.05901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.497001  V
** inner: 0.679001  V


.END