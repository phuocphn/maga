** Name: two_stage_single_output_op_amp_79_5

.MACRO two_stage_single_output_op_amp_79_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=13e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=7e-6 W=141e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=354e-6
mMainBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=166e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=31e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mFoldedCascodeFirstStageLoad10 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=10e-6 W=86e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=22e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=22e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=123e-6
mMainBias14 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=269e-6
mSecondStage1Transconductor15 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=195e-6
mFoldedCascodeFirstStageLoad16 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=86e-6
mMainBias17 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=51e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=25e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=23e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=23e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=354e-6
mFoldedCascodeFirstStageLoad23 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=25e-6
mMainBias24 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=26e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_79_5

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 8.82201 mW
** Area: 10395 (mu_m)^2
** Transit frequency: 5.07401 MHz
** Transit frequency with error factor: 5.07398 MHz
** Slew rate: 3.5451 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 3.49001 V
** VoutMin: 0.410001 V
** VcmMax: 4.71001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorNmos: 3.94161e+07 muA
** NormalTransistorNmos: 2.04518e+08 muA
** NormalTransistorPmos: -3.24769e+07 muA
** NormalTransistorPmos: -1.64489e+07 muA
** NormalTransistorPmos: -2.81999e+07 muA
** NormalTransistorPmos: -1.64469e+07 muA
** NormalTransistorPmos: -2.81979e+07 muA
** NormalTransistorNmos: 1.64481e+07 muA
** NormalTransistorNmos: 1.64471e+07 muA
** NormalTransistorNmos: 1.64461e+07 muA
** NormalTransistorNmos: 1.64471e+07 muA
** NormalTransistorNmos: 2.35001e+07 muA
** NormalTransistorNmos: 2.35011e+07 muA
** NormalTransistorNmos: 1.17501e+07 muA
** NormalTransistorNmos: 1.17501e+07 muA
** NormalTransistorNmos: 1.42152e+09 muA
** NormalTransistorPmos: -1.42151e+09 muA
** DiodeTransistorPmos: -1.42151e+09 muA
** DiodeTransistorNmos: 3.24761e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.94169e+07 muA
** NormalTransistorPmos: -3.94179e+07 muA
** DiodeTransistorPmos: -2.04517e+08 muA
** DiodeTransistorPmos: -2.04518e+08 muA


** Expected Voltages: 
** ibias: 0.674001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.42601  V
** out: 2.5  V
** outFirstStage: 0.819001  V
** outInputVoltageBiasXXpXX1: 2.92401  V
** outSourceVoltageBiasXXpXX1: 3.96401  V
** outSourceVoltageBiasXXpXX2: 3.74001  V
** outVoltageBiasXXnXX1: 1.02401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.469001  V
** innerTransistorStack1Load2: 0.468001  V
** innerTransistorStack2Load2: 0.468001  V
** out1: 0.619001  V
** sourceGCC1: 3.49601  V
** sourceGCC2: 3.49601  V
** sourceTransconductance: 1.93601  V
** inner: 3.95601  V


.END