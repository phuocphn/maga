** Name: two_stage_single_output_op_amp_54_5

.MACRO two_stage_single_output_op_amp_54_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mMainBias3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=4e-6 W=125e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=6e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=552e-6
mMainBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=124e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=87e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=120e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=120e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=80e-6
mMainBias13 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=317e-6
mSecondStage1Transconductor14 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=296e-6
mFoldedCascodeFirstStageLoad15 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=87e-6
mMainBias16 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=569e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=38e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=38e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=6e-6
mMainBias21 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=26e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=552e-6
mFoldedCascodeFirstStageLoad23 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=569e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.2001e-12
.EOM two_stage_single_output_op_amp_54_5

** Expected Performance Values: 
** Gain: 135 dB
** Power consumption: 9.40301 mW
** Area: 13578 (mu_m)^2
** Transit frequency: 3.88701 MHz
** Transit frequency with error factor: 3.88747 MHz
** Slew rate: 3.50022 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 3 V
** VoutMin: 0.320001 V
** VcmMax: 4.66001 V
** VcmMin: 0.75 V


** Expected Currents: 
** NormalTransistorNmos: 1.37341e+07 muA
** NormalTransistorNmos: 3.14756e+08 muA
** NormalTransistorPmos: -6.50579e+07 muA
** NormalTransistorPmos: -5.72189e+07 muA
** NormalTransistorPmos: -9.64569e+07 muA
** NormalTransistorPmos: -5.72189e+07 muA
** NormalTransistorPmos: -9.64569e+07 muA
** NormalTransistorNmos: 5.72181e+07 muA
** NormalTransistorNmos: 5.72171e+07 muA
** NormalTransistorNmos: 5.72181e+07 muA
** NormalTransistorNmos: 5.72171e+07 muA
** NormalTransistorNmos: 7.84791e+07 muA
** NormalTransistorNmos: 3.92391e+07 muA
** NormalTransistorNmos: 3.92391e+07 muA
** NormalTransistorNmos: 1.28416e+09 muA
** NormalTransistorPmos: -1.28415e+09 muA
** DiodeTransistorPmos: -1.28415e+09 muA
** DiodeTransistorNmos: 6.50571e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.37349e+07 muA
** NormalTransistorPmos: -1.37359e+07 muA
** DiodeTransistorPmos: -3.14755e+08 muA
** DiodeTransistorPmos: -3.14754e+08 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.931001  V
** inputVoltageBiasXXpXX2: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.726001  V
** outInputVoltageBiasXXpXX1: 2.43601  V
** outSourceVoltageBiasXXpXX1: 3.71801  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.89801  V
** inner: 3.71301  V


.END