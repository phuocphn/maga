** Name: two_stage_single_output_op_amp_6_2

.MACRO two_stage_single_output_op_amp_6_2 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=25e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=6e-6 W=25e-6
mSecondStage1StageBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=27e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=12e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=6e-6 W=25e-6
mSecondStage1Transconductor6 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=124e-6
mSecondStage1Transconductor7 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=351e-6
mSimpleFirstStageLoad8 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=25e-6
mSimpleFirstStageTransconductor9 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=16e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=79e-6
mSecondStage1StageBias11 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=426e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=16e-6
mMainBias13 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=254e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_6_2

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 3.27501 mW
** Area: 5977 (mu_m)^2
** Transit frequency: 3.16601 MHz
** Transit frequency with error factor: 3.15509 MHz
** Slew rate: 13.6014 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** negPSRR: 90 dB
** posPSRR: 98 dB
** VoutMax: 4.63001 V
** VoutMin: 0.75 V
** VcmMax: 3.38001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorPmos: -2.14912e+08 muA
** DiodeTransistorNmos: 3.34211e+07 muA
** NormalTransistorNmos: 3.34201e+07 muA
** NormalTransistorNmos: 3.34211e+07 muA
** DiodeTransistorNmos: 3.34201e+07 muA
** NormalTransistorPmos: -6.68429e+07 muA
** NormalTransistorPmos: -3.34219e+07 muA
** NormalTransistorPmos: -3.34219e+07 muA
** NormalTransistorNmos: 3.53309e+08 muA
** NormalTransistorNmos: 3.53308e+08 muA
** NormalTransistorPmos: -3.53308e+08 muA
** DiodeTransistorNmos: 2.14913e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.06101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.889001  V
** outVoltageBiasXXnXX1: 1.15501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 1.29401  V
** innerTransistorStack1Load1: 0.711001  V
** innerTransistorStack2Load1: 0.712001  V
** sourceTransconductance: 3.74501  V
** innerTransconductance: 0.484001  V


.END