** Name: two_stage_single_output_op_amp_78_6

.MACRO two_stage_single_output_op_amp_78_6 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=108e-6
mFoldedCascodeFirstStageLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=2e-6 W=93e-6
mMainBias3 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=40e-6
mSecondStage1StageBias4 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=433e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=5e-6
mMainBias7 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=563e-6
mMainBias9 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=2e-6 W=93e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=64e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=64e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=433e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=38e-6
mMainBias15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=40e-6
mSecondStage1Transconductor16 out inputVoltageBiasXXnXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=437e-6
mFoldedCascodeFirstStageLoad17 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=108e-6
mMainBias18 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=29e-6
mMainBias19 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=174e-6
mFoldedCascodeFirstStageLoad20 FirstStageYinnerOutputLoad2 outInputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=103e-6
mFoldedCascodeFirstStageLoad21 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=162e-6
mFoldedCascodeFirstStageLoad22 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=162e-6
mMainBias23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias24 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=381e-6
mSecondStage1StageBias25 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=563e-6
mFoldedCascodeFirstStageLoad26 outFirstStage outInputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=103e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.1001e-12
.EOM two_stage_single_output_op_amp_78_6

** Expected Performance Values: 
** Gain: 164 dB
** Power consumption: 7.86001 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 3.81201 MHz
** Transit frequency with error factor: 3.81175 MHz
** Slew rate: 7.26206 V/mu_s
** Phase margin: 66.4632°
** CMRR: 139 dB
** VoutMax: 3.62001 V
** VoutMin: 0.660001 V
** VcmMax: 5.17001 V
** VcmMin: 1.43001 V


** Expected Currents: 
** NormalTransistorNmos: 7.25401e+06 muA
** NormalTransistorNmos: 4.35341e+07 muA
** NormalTransistorPmos: -3.66975e+08 muA
** NormalTransistorPmos: -1.0285e+08 muA
** NormalTransistorPmos: -1.55946e+08 muA
** NormalTransistorPmos: -1.0285e+08 muA
** NormalTransistorPmos: -1.55946e+08 muA
** DiodeTransistorNmos: 1.02851e+08 muA
** DiodeTransistorNmos: 1.0285e+08 muA
** NormalTransistorNmos: 1.02851e+08 muA
** NormalTransistorNmos: 1.0285e+08 muA
** NormalTransistorNmos: 1.06191e+08 muA
** DiodeTransistorNmos: 1.06192e+08 muA
** NormalTransistorNmos: 5.30951e+07 muA
** NormalTransistorNmos: 5.30951e+07 muA
** NormalTransistorNmos: 8.32323e+08 muA
** NormalTransistorNmos: 8.32322e+08 muA
** NormalTransistorPmos: -8.32322e+08 muA
** DiodeTransistorPmos: -8.32323e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 3.66976e+08 muA
** DiodeTransistorPmos: -7.25499e+06 muA
** NormalTransistorPmos: -7.25599e+06 muA
** DiodeTransistorPmos: -4.35349e+07 muA
** DiodeTransistorPmos: -4.35359e+07 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.06601  V
** out: 2.5  V
** outFirstStage: 0.916001  V
** outInputVoltageBiasXXpXX1: 3.05901  V
** outInputVoltageBiasXXpXX2: 3.14501  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.03101  V
** outSourceVoltageBiasXXpXX2: 4.20501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 1.12101  V
** innerTransistorStack1Load2: 0.566001  V
** innerTransistorStack2Load2: 0.566001  V
** sourceGCC1: 3.94501  V
** sourceGCC2: 3.94501  V
** sourceTransconductance: 1.78101  V
** innerTransconductance: 0.511001  V
** inner: 0.556001  V
** inner: 4.02401  V


.END