** Name: symmetrical_op_amp25

.MACRO symmetrical_op_amp25 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=11e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSecondStage1StageBias3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=78e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=16e-6
mSymmetricalFirstStageLoad6 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=78e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=258e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias9 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=258e-6
mMainBias10 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos4 L=5e-6 W=112e-6
mSymmetricalFirstStageTransconductor11 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=105e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias12 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=3e-6 W=96e-6
mMainBias13 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=12e-6
mSecondStage1StageBias14 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=96e-6
mSymmetricalFirstStageTransconductor15 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=105e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=85e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=85e-6
mMainBias18 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=48e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor19 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=199e-6
mSecondStage1Transconductor20 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=199e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp25

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 6.55001 mW
** Area: 7413 (mu_m)^2
** Transit frequency: 19.0701 MHz
** Transit frequency with error factor: 19.0703 MHz
** Slew rate: 30.2875 V/mu_s
** Phase margin: 81.933°
** CMRR: 137 dB
** negPSRR: 60 dB
** posPSRR: 52 dB
** VoutMax: 4.26001 V
** VoutMin: 0.540001 V
** VcmMax: 4.40001 V
** VcmMin: 0.880001 V


** Expected Currents: 
** NormalTransistorNmos: 1.09501e+07 muA
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -3.23469e+07 muA
** DiodeTransistorPmos: -2.73758e+08 muA
** DiodeTransistorPmos: -2.73758e+08 muA
** NormalTransistorNmos: 5.47516e+08 muA
** NormalTransistorNmos: 2.73759e+08 muA
** NormalTransistorNmos: 2.73759e+08 muA
** NormalTransistorNmos: 3.03829e+08 muA
** NormalTransistorNmos: 3.03828e+08 muA
** NormalTransistorPmos: -3.03828e+08 muA
** NormalTransistorPmos: -3.03827e+08 muA
** NormalTransistorNmos: 3.03829e+08 muA
** NormalTransistorNmos: 3.03828e+08 muA
** NormalTransistorPmos: -3.03828e+08 muA
** NormalTransistorPmos: -3.03827e+08 muA
** DiodeTransistorNmos: 3.23461e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.09509e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 0.636001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.943001  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 3.99101  V
** innerComplementarySecondStage: 0.609001  V
** inputVoltageBiasXXpXX0: 3.92001  V
** out: 2.5  V
** outFirstStage: 3.99101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.84601  V
** innerStageBias: 0.204001  V
** innerTransconductance: 4.54101  V
** inner: 0.204001  V
** inner: 4.54101  V


.END