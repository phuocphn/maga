** Name: two_stage_single_output_op_amp_36_7

.MACRO two_stage_single_output_op_amp_36_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=9e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=14e-6
mSimpleFirstStageLoad4 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=9e-6 W=63e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=212e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=16e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=17e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=14e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mMainBias10 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=348e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=17e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=212e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=297e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=9e-6 W=63e-6
mMainBias16 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=39e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_36_7

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 2.38401 mW
** Area: 8973 (mu_m)^2
** Transit frequency: 2.60101 MHz
** Transit frequency with error factor: 2.59794 MHz
** Slew rate: 4.19552 V/mu_s
** Phase margin: 61.8795°
** CMRR: 100 dB
** negPSRR: 95 dB
** posPSRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 0.210001 V
** VcmMax: 3.85001 V
** VcmMin: 1.82001 V


** Expected Currents: 
** NormalTransistorNmos: 4.92901e+06 muA
** NormalTransistorPmos: -1.21769e+07 muA
** DiodeTransistorPmos: -9.48599e+06 muA
** DiodeTransistorPmos: -9.48699e+06 muA
** NormalTransistorPmos: -9.48799e+06 muA
** NormalTransistorPmos: -9.48699e+06 muA
** NormalTransistorNmos: 1.89731e+07 muA
** DiodeTransistorNmos: 1.89721e+07 muA
** NormalTransistorNmos: 9.48701e+06 muA
** NormalTransistorNmos: 9.48701e+06 muA
** NormalTransistorNmos: 4.30794e+08 muA
** NormalTransistorPmos: -4.30793e+08 muA
** DiodeTransistorNmos: 1.21761e+07 muA
** NormalTransistorNmos: 1.21751e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.92999e+06 muA


** Expected Voltages: 
** ibias: 0.615001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.25  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.56601  V
** outSourceVoltageBiasXXnXX1: 0.783001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.44801  V
** innerSourceLoad1: 4.28601  V
** innerTransistorStack2Load1: 4.28701  V
** sourceTransconductance: 1.83701  V
** inner: 0.780001  V


.END