** Name: two_stage_single_output_op_amp_5_5

.MACRO two_stage_single_output_op_amp_5_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=42e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=22e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=341e-6
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=257e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=110e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=110e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=535e-6
mSimpleFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=257e-6
mMainBias11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=10e-6
mSimpleFirstStageTransconductor12 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=107e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=581e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=32e-6
mSecondStage1StageBias16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=341e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=107e-6
mMainBias18 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=227e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_5_5

** Expected Performance Values: 
** Gain: 106 dB
** Power consumption: 6.53901 mW
** Area: 9436 (mu_m)^2
** Transit frequency: 25.1861 MHz
** Transit frequency with error factor: 25.1658 MHz
** Slew rate: 30.2678 V/mu_s
** Phase margin: 66.4632°
** CMRR: 104 dB
** negPSRR: 106 dB
** posPSRR: 234 dB
** VoutMax: 3.61001 V
** VoutMin: 0.150001 V
** VcmMax: 4.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 6.70801e+07 muA
** NormalTransistorPmos: -5.38019e+07 muA
** NormalTransistorPmos: -7.69599e+06 muA
** NormalTransistorNmos: 6.99531e+07 muA
** NormalTransistorNmos: 6.99521e+07 muA
** NormalTransistorNmos: 6.99511e+07 muA
** NormalTransistorNmos: 6.99521e+07 muA
** NormalTransistorPmos: -1.39902e+08 muA
** NormalTransistorPmos: -6.99519e+07 muA
** NormalTransistorPmos: -6.99519e+07 muA
** NormalTransistorNmos: 1.01931e+09 muA
** NormalTransistorPmos: -1.0193e+09 muA
** DiodeTransistorPmos: -1.01931e+09 muA
** DiodeTransistorNmos: 5.38011e+07 muA
** DiodeTransistorNmos: 7.69501e+06 muA
** DiodeTransistorPmos: -6.70809e+07 muA
** NormalTransistorPmos: -6.70799e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.20501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.05001  V
** outSourceVoltageBiasXXpXX1: 4.02501  V
** outVoltageBiasXXnXX0: 1.14701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.25501  V
** inner: 4.02601  V


.END