** Name: two_stage_single_output_op_amp_20_1

.MACRO two_stage_single_output_op_amp_20_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=65e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=12e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=107e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=65e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=496e-6
mSimpleFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=10e-6 W=12e-6
mMainBias10 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSimpleFirstStageTransconductor11 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=129e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=107e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=12e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mSecondStage1StageBias15 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=190e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=129e-6
mMainBias17 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_20_1

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 1.17801 mW
** Area: 7317 (mu_m)^2
** Transit frequency: 4.48801 MHz
** Transit frequency with error factor: 4.48382 MHz
** Slew rate: 5.46811 V/mu_s
** Phase margin: 63.5984°
** CMRR: 104 dB
** negPSRR: 106 dB
** posPSRR: 156 dB
** VoutMax: 4.78001 V
** VoutMin: 0.150001 V
** VcmMax: 3.28001 V
** VcmMin: 0.340001 V


** Expected Currents: 
** NormalTransistorNmos: 2.82801e+06 muA
** NormalTransistorPmos: -8.49899e+06 muA
** NormalTransistorPmos: -2.12059e+07 muA
** DiodeTransistorNmos: 1.23811e+07 muA
** NormalTransistorNmos: 1.23811e+07 muA
** NormalTransistorNmos: 1.23811e+07 muA
** NormalTransistorPmos: -2.47649e+07 muA
** DiodeTransistorPmos: -2.47659e+07 muA
** NormalTransistorPmos: -1.23819e+07 muA
** NormalTransistorPmos: -1.23819e+07 muA
** NormalTransistorNmos: 1.58299e+08 muA
** NormalTransistorPmos: -1.58298e+08 muA
** DiodeTransistorNmos: 8.49801e+06 muA
** DiodeTransistorNmos: 2.12051e+07 muA
** DiodeTransistorPmos: -2.82899e+06 muA
** NormalTransistorPmos: -2.82999e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.903001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.47601  V
** outSourceVoltageBiasXXpXX1: 4.23801  V
** outVoltageBiasXXnXX0: 0.588001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.25701  V
** inner: 4.23801  V


.END