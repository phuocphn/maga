** Name: two_stage_single_output_op_amp_130_6

.MACRO two_stage_single_output_op_amp_130_6 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=116e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=71e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=45e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=124e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=145e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=145e-6
mSimpleFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=486e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=212e-6
mMainBias11 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=71e-6
mSecondStage1Transconductor12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=524e-6
mSimpleFirstStageLoad13 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=486e-6
mSimpleFirstStageTransconductor14 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=95e-6
mSimpleFirstStageLoad15 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=71e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=305e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=45e-6
mMainBias18 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=290e-6
mSecondStage1StageBias19 out inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=124e-6
mSimpleFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=6e-6 W=108e-6
mSimpleFirstStageTransconductor21 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=95e-6
mMainBias22 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=27e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.4001e-12
.EOM two_stage_single_output_op_amp_130_6

** Expected Performance Values: 
** Gain: 135 dB
** Power consumption: 7.27401 mW
** Area: 9353 (mu_m)^2
** Transit frequency: 4.45501 MHz
** Transit frequency with error factor: 4.44733 MHz
** Slew rate: 12.4067 V/mu_s
** Phase margin: 60.1606°
** CMRR: 82 dB
** VoutMax: 3.58001 V
** VoutMin: 0.310001 V
** VcmMax: 3.40001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 1.48553e+08 muA
** NormalTransistorPmos: -2.2625e+07 muA
** NormalTransistorPmos: -2.42705e+08 muA
** NormalTransistorPmos: -1.79674e+08 muA
** NormalTransistorPmos: -1.79674e+08 muA
** DiodeTransistorPmos: -1.79674e+08 muA
** NormalTransistorNmos: 3.08551e+08 muA
** NormalTransistorNmos: 3.0855e+08 muA
** NormalTransistorNmos: 3.08551e+08 muA
** NormalTransistorNmos: 3.0855e+08 muA
** NormalTransistorPmos: -2.5775e+08 muA
** NormalTransistorPmos: -1.28875e+08 muA
** NormalTransistorPmos: -1.28875e+08 muA
** NormalTransistorNmos: 4.03781e+08 muA
** NormalTransistorNmos: 4.03782e+08 muA
** NormalTransistorPmos: -4.0378e+08 muA
** DiodeTransistorPmos: -4.03781e+08 muA
** DiodeTransistorNmos: 2.26241e+07 muA
** DiodeTransistorNmos: 2.42706e+08 muA
** DiodeTransistorPmos: -1.48552e+08 muA
** NormalTransistorPmos: -1.48553e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.563001  V
** inputVoltageBiasXXpXX1: 3.01401  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.00701  V
** outVoltageBiasXXnXX1: 0.720001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.165001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.165001  V
** out1: 2.37201  V
** sourceTransconductance: 3.79001  V
** innerTransconductance: 0.150001  V
** inner: 4.00601  V


.END