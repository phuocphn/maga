** Name: symmetrical_op_amp191

.MACRO symmetrical_op_amp191 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=12e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=96e-6
mSymmetricalFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=129e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=36e-6
mMainBias5 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=12e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=129e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=96e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mSymmetricalFirstStageTransconductor10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=14e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=18e-6
mSymmetricalFirstStageTransconductor12 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=14e-6
mMainBias13 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=123e-6
mMainBias14 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=14e-6
mSymmetricalFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=74e-6
mSymmetricalFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=73e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=87e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=87e-6
mSymmetricalFirstStageLoad19 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=131e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor20 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=156e-6
mSecondStage1Transconductor21 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=156e-6
mSymmetricalFirstStageLoad22 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=131e-6
mMainBias23 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=266e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp191

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 3.04001 mW
** Area: 6854 (mu_m)^2
** Transit frequency: 4.66701 MHz
** Transit frequency with error factor: 4.66706 MHz
** Slew rate: 6.26986 V/mu_s
** Phase margin: 74.4846°
** CMRR: 137 dB
** negPSRR: 129 dB
** posPSRR: 62 dB
** VoutMax: 4.25 V
** VoutMin: 0.580001 V
** VcmMax: 4.81001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 1.16571e+07 muA
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -2.5375e+08 muA
** NormalTransistorPmos: -5.26909e+07 muA
** NormalTransistorPmos: -5.26919e+07 muA
** NormalTransistorPmos: -5.26909e+07 muA
** NormalTransistorPmos: -5.26919e+07 muA
** NormalTransistorNmos: 1.05382e+08 muA
** DiodeTransistorNmos: 1.05383e+08 muA
** NormalTransistorNmos: 5.26901e+07 muA
** NormalTransistorNmos: 5.26901e+07 muA
** NormalTransistorNmos: 6.28151e+07 muA
** NormalTransistorNmos: 6.28141e+07 muA
** NormalTransistorPmos: -6.28159e+07 muA
** NormalTransistorPmos: -6.28149e+07 muA
** DiodeTransistorNmos: 6.28151e+07 muA
** NormalTransistorPmos: -6.28159e+07 muA
** NormalTransistorPmos: -6.28149e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 2.5375e+08 muA
** DiodeTransistorPmos: -1.16579e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 1.15101  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.580001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.576001  V
** outVoltageBiasXXnXX2: 0.985001  V
** outVoltageBiasXXpXX0: 3.97201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.88401  V
** innerStageBias: 0.175001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V
** inner: 0.574001  V


.END