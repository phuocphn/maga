** Name: two_stage_single_output_op_amp_50_7

.MACRO two_stage_single_output_op_amp_50_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=69e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=115e-6
mFoldedCascodeFirstStageTransconductor5 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=33e-6
mFoldedCascodeFirstStageTransconductor6 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=33e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=12e-6
mSecondStage1StageBias8 out ibias sourceNmos sourceNmos nmos4 L=7e-6 W=507e-6
mFoldedCascodeFirstStageLoad9 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
mMainBias10 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=47e-6
mFoldedCascodeFirstStageLoad11 FirstStageYout1 outInputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageLoad12 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=210e-6
mFoldedCascodeFirstStageLoad15 outFirstStage outInputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=16e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_50_7

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 4.18801 mW
** Area: 5769 (mu_m)^2
** Transit frequency: 3.60501 MHz
** Transit frequency with error factor: 3.60113 MHz
** Slew rate: 3.72734 V/mu_s
** Phase margin: 65.3172°
** CMRR: 106 dB
** VoutMax: 4.25 V
** VoutMin: 0.340001 V
** VcmMax: 5.23001 V
** VcmMin: 0.910001 V


** Expected Currents: 
** NormalTransistorNmos: 6.65081e+07 muA
** NormalTransistorPmos: -1.68069e+07 muA
** NormalTransistorPmos: -2.52089e+07 muA
** NormalTransistorPmos: -1.68089e+07 muA
** NormalTransistorPmos: -2.52129e+07 muA
** DiodeTransistorNmos: 1.68081e+07 muA
** NormalTransistorNmos: 1.68081e+07 muA
** NormalTransistorNmos: 1.68061e+07 muA
** NormalTransistorNmos: 8.40301e+06 muA
** NormalTransistorNmos: 8.40301e+06 muA
** NormalTransistorNmos: 7.10738e+08 muA
** NormalTransistorPmos: -7.10737e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.65089e+07 muA
** DiodeTransistorPmos: -6.65099e+07 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXpXX1: 3.46001  V
** outSourceVoltageBiasXXpXX1: 4.25701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.612001  V
** sourceGCC1: 4.26601  V
** sourceGCC2: 4.26601  V
** sourceTransconductance: 1.93001  V


.END