** Name: two_stage_single_output_op_amp_29_10

.MACRO two_stage_single_output_op_amp_29_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=310e-6
mMainBias4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=89e-6
mSecondStage1StageBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=300e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=36e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=158e-6
mMainBias9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
mMainBias10 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=66e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=36e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSecondStage1Transconductor14 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=310e-6
mMainBias16 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=530e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.7001e-12
.EOM two_stage_single_output_op_amp_29_10

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 8.90601 mW
** Area: 7571 (mu_m)^2
** Transit frequency: 9.68001 MHz
** Transit frequency with error factor: 9.62475 MHz
** Slew rate: 32.437 V/mu_s
** Phase margin: 60.1606°
** CMRR: 83 dB
** negPSRR: 115 dB
** posPSRR: 81 dB
** VoutMax: 4.39001 V
** VoutMin: 0.200001 V
** VcmMax: 4.54001 V
** VcmMin: 1.95001 V


** Expected Currents: 
** NormalTransistorNmos: 2.30011e+07 muA
** NormalTransistorNmos: 1.10621e+08 muA
** NormalTransistorPmos: -1.3891e+08 muA
** DiodeTransistorPmos: -2.47295e+08 muA
** NormalTransistorPmos: -2.47295e+08 muA
** NormalTransistorNmos: 4.9459e+08 muA
** NormalTransistorNmos: 4.94589e+08 muA
** NormalTransistorNmos: 2.47296e+08 muA
** NormalTransistorNmos: 2.47296e+08 muA
** NormalTransistorNmos: 1.00409e+09 muA
** NormalTransistorPmos: -1.00408e+09 muA
** NormalTransistorPmos: -1.00408e+09 muA
** DiodeTransistorNmos: 1.38911e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.30019e+07 muA
** DiodeTransistorPmos: -1.1062e+08 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.19501  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.13101  V
** outVoltageBiasXXnXX1: 0.809001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.211001  V
** out1: 4.13601  V
** sourceTransconductance: 1.34501  V
** innerTransconductance: 4.55501  V


.END