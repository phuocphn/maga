** Name: symmetrical_op_amp7

.MACRO symmetrical_op_amp7 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=125e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=13e-6
mSymmetricalFirstStageLoad4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=125e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=90e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=5e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=182e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=182e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=4e-6 W=30e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=30e-6
mMainBias12 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=13e-6
mSymmetricalFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=158e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=90e-6
mMainBias15 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mSymmetricalFirstStageTransconductor16 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=115e-6
mMainBias17 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=126e-6
mSymmetricalFirstStageTransconductor19 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=115e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 2.36801 mW
** Area: 5188 (mu_m)^2
** Transit frequency: 3.12901 MHz
** Transit frequency with error factor: 3.12878 MHz
** Slew rate: 11.5362 V/mu_s
** Phase margin: 84.7978°
** CMRR: 135 dB
** negPSRR: 34 dB
** posPSRR: 36 dB
** VoutMax: 4.34001 V
** VoutMin: 0.570001 V
** VcmMax: 3.61001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 1.69211e+07 muA
** NormalTransistorPmos: -1.71839e+07 muA
** NormalTransistorPmos: -2.82709e+07 muA
** DiodeTransistorNmos: 8.00951e+07 muA
** DiodeTransistorNmos: 8.00951e+07 muA
** NormalTransistorPmos: -1.60191e+08 muA
** NormalTransistorPmos: -8.00959e+07 muA
** NormalTransistorPmos: -8.00959e+07 muA
** NormalTransistorNmos: 1.15548e+08 muA
** NormalTransistorNmos: 1.15549e+08 muA
** NormalTransistorPmos: -1.15547e+08 muA
** NormalTransistorPmos: -1.15548e+08 muA
** DiodeTransistorPmos: -1.15547e+08 muA
** NormalTransistorNmos: 1.15548e+08 muA
** NormalTransistorNmos: 1.15549e+08 muA
** DiodeTransistorNmos: 1.71831e+07 muA
** DiodeTransistorNmos: 2.82701e+07 muA
** DiodeTransistorPmos: -1.69219e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.980001  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 4.16701  V
** inputVoltageBiasXXnXX0: 0.778001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.65401  V
** innerStageBias: 4.64101  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END