** Name: two_stage_single_output_op_amp_205_10

.MACRO two_stage_single_output_op_amp_205_10 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=20e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=20e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias4 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=158e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=78e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=45e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=20e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=174e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=132e-6
mMainBias11 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=59e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=508e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=2e-6 W=20e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=174e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=316e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=325e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=325e-6
mSimpleFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=569e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=424e-6
mMainBias20 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=160e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=569e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.2001e-12
.EOM two_stage_single_output_op_amp_205_10

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 14.7491 mW
** Area: 12600 (mu_m)^2
** Transit frequency: 6.72901 MHz
** Transit frequency with error factor: 6.72546 MHz
** Slew rate: 6.34163 V/mu_s
** Phase margin: 60.1606°
** CMRR: 111 dB
** VoutMax: 4.25 V
** VoutMin: 0.340001 V
** VcmMax: 4.78001 V
** VcmMin: 1.47001 V


** Expected Currents: 
** NormalTransistorNmos: 7.9008e+08 muA
** NormalTransistorNmos: 1.44595e+08 muA
** NormalTransistorPmos: -1.48164e+08 muA
** DiodeTransistorNmos: 2.3989e+08 muA
** NormalTransistorNmos: 2.39891e+08 muA
** NormalTransistorNmos: 2.39892e+08 muA
** DiodeTransistorNmos: 2.39891e+08 muA
** NormalTransistorPmos: -2.95124e+08 muA
** NormalTransistorPmos: -2.95125e+08 muA
** NormalTransistorPmos: -2.95126e+08 muA
** NormalTransistorPmos: -2.95125e+08 muA
** NormalTransistorNmos: 1.1047e+08 muA
** NormalTransistorNmos: 1.10469e+08 muA
** NormalTransistorNmos: 5.52351e+07 muA
** NormalTransistorNmos: 5.52351e+07 muA
** NormalTransistorNmos: 1.26676e+09 muA
** NormalTransistorPmos: -1.26675e+09 muA
** NormalTransistorPmos: -1.26675e+09 muA
** DiodeTransistorNmos: 1.48165e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.90079e+08 muA
** DiodeTransistorPmos: -1.44594e+08 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.06401  V
** inputVoltageBiasXXpXX2: 3.98301  V
** out: 2.5  V
** outFirstStage: 4.02801  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.486001  V
** innerTransistorStack1Load1: 1.15601  V
** innerTransistorStack1Load2: 4.42001  V
** innerTransistorStack2Load2: 4.42001  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.59201  V


.END