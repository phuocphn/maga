** Name: two_stage_single_output_op_amp_16_2

.MACRO two_stage_single_output_op_amp_16_2 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=27e-6
mSecondStage1StageBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=130e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=23e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=317e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=60e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=385e-6
mSecondStage1Transconductor8 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=169e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=27e-6
mMainBias10 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=306e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=60e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=317e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=110e-6
mSecondStage1StageBias15 out ibias sourcePmos sourcePmos pmos4 L=5e-6 W=402e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mMainBias17 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=80e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_16_2

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 1.90201 mW
** Area: 14818 (mu_m)^2
** Transit frequency: 2.65001 MHz
** Transit frequency with error factor: 2.64696 MHz
** Slew rate: 3.50004 V/mu_s
** Phase margin: 71.6198°
** CMRR: 96 dB
** negPSRR: 98 dB
** posPSRR: 125 dB
** VoutMax: 4.65001 V
** VoutMin: 0.370001 V
** VcmMax: 3.02001 V
** VcmMin: 0.0300001 V


** Expected Currents: 
** NormalTransistorNmos: 8.32601e+07 muA
** NormalTransistorPmos: -3.53779e+07 muA
** NormalTransistorPmos: -4.80969e+07 muA
** DiodeTransistorNmos: 7.89401e+06 muA
** NormalTransistorNmos: 7.89401e+06 muA
** NormalTransistorPmos: -1.57909e+07 muA
** DiodeTransistorPmos: -1.57919e+07 muA
** NormalTransistorPmos: -7.89499e+06 muA
** NormalTransistorPmos: -7.89499e+06 muA
** NormalTransistorNmos: 1.77779e+08 muA
** NormalTransistorNmos: 1.77778e+08 muA
** NormalTransistorPmos: -1.77778e+08 muA
** DiodeTransistorNmos: 3.53771e+07 muA
** DiodeTransistorNmos: 4.80961e+07 muA
** DiodeTransistorPmos: -8.32609e+07 muA
** NormalTransistorPmos: -8.32619e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.08601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.780001  V
** out: 2.5  V
** outFirstStage: 0.586001  V
** outInputVoltageBiasXXpXX1: 3.22801  V
** outSourceVoltageBiasXXpXX1: 4.11401  V
** outVoltageBiasXXnXX0: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.590001  V
** sourceTransconductance: 3.27401  V
** innerTransconductance: 0.181001  V
** inner: 4.11201  V


.END