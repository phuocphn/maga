** Name: two_stage_single_output_op_amp_189_12

.MACRO two_stage_single_output_op_amp_189_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=8e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=13e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=283e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=34e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=179e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=187e-6
mSimpleFirstStageLoad10 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=71e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=283e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=1e-6 W=21e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=187e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=150e-6
mMainBias17 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=61e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=555e-6
mSimpleFirstStageLoad19 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=555e-6
mSimpleFirstStageLoad20 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=496e-6
mSecondStage1Transconductor21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=564e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
mSimpleFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=496e-6
mMainBias24 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=55e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.7001e-12
.EOM two_stage_single_output_op_amp_189_12

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 14.9991 mW
** Area: 10082 (mu_m)^2
** Transit frequency: 10.5891 MHz
** Transit frequency with error factor: 10.583 MHz
** Slew rate: 9.97969 V/mu_s
** Phase margin: 60.1606°
** CMRR: 117 dB
** VoutMax: 4.25 V
** VoutMin: 1.26001 V
** VcmMax: 4.77001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 9.95231e+07 muA
** NormalTransistorNmos: 4.03661e+07 muA
** NormalTransistorPmos: -6.64939e+07 muA
** NormalTransistorNmos: 6.00276e+08 muA
** NormalTransistorNmos: 6.00277e+08 muA
** DiodeTransistorNmos: 6.00276e+08 muA
** NormalTransistorPmos: -6.59636e+08 muA
** NormalTransistorPmos: -6.59637e+08 muA
** NormalTransistorPmos: -6.59637e+08 muA
** NormalTransistorPmos: -6.59637e+08 muA
** NormalTransistorNmos: 1.18722e+08 muA
** NormalTransistorNmos: 1.18721e+08 muA
** NormalTransistorNmos: 5.93611e+07 muA
** NormalTransistorNmos: 5.93611e+07 muA
** NormalTransistorNmos: 1.46424e+09 muA
** DiodeTransistorNmos: 1.46424e+09 muA
** NormalTransistorPmos: -1.46423e+09 muA
** NormalTransistorPmos: -1.46423e+09 muA
** DiodeTransistorNmos: 6.64931e+07 muA
** NormalTransistorNmos: 6.64921e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.95239e+07 muA
** DiodeTransistorPmos: -4.03669e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.05401  V
** outInputVoltageBiasXXnXX1: 1.66401  V
** outSourceVoltageBiasXXnXX1: 0.832001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.07001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.14701  V
** innerStageBias: 0.524001  V
** innerTransistorStack1Load2: 4.52201  V
** innerTransistorStack2Load2: 4.52201  V
** out1: 2.13601  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.61801  V
** inner: 0.832001  V


.END