** Name: two_stage_single_output_op_amp_73_10

.MACRO two_stage_single_output_op_amp_73_10 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=33e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=118e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=46e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=119e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=119e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=414e-6
mMainBias11 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=57e-6
mMainBias12 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=26e-6
mSecondStage1StageBias13 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=534e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=5e-6 W=101e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=201e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=257e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=257e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=472e-6
mSecondStage1Transconductor19 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=201e-6
mMainBias21 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=347e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.5e-12
.EOM two_stage_single_output_op_amp_73_10

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 10.0801 mW
** Area: 9743 (mu_m)^2
** Transit frequency: 6.83901 MHz
** Transit frequency with error factor: 6.83897 MHz
** Slew rate: 4.64303 V/mu_s
** Phase margin: 60.1606°
** CMRR: 144 dB
** VoutMax: 4.25 V
** VoutMin: 0.340001 V
** VcmMax: 5.23001 V
** VcmMin: 1.45001 V


** Expected Currents: 
** NormalTransistorNmos: 1.42147e+08 muA
** NormalTransistorNmos: 6.37201e+07 muA
** NormalTransistorPmos: -1.89206e+08 muA
** NormalTransistorPmos: -8.16329e+07 muA
** NormalTransistorPmos: -1.38296e+08 muA
** NormalTransistorPmos: -8.16329e+07 muA
** NormalTransistorPmos: -1.38296e+08 muA
** NormalTransistorNmos: 8.16321e+07 muA
** NormalTransistorNmos: 8.16321e+07 muA
** DiodeTransistorNmos: 8.16321e+07 muA
** NormalTransistorNmos: 1.13326e+08 muA
** NormalTransistorNmos: 1.13325e+08 muA
** NormalTransistorNmos: 5.66631e+07 muA
** NormalTransistorNmos: 5.66631e+07 muA
** NormalTransistorNmos: 1.33431e+09 muA
** NormalTransistorPmos: -1.3343e+09 muA
** NormalTransistorPmos: -1.3343e+09 muA
** DiodeTransistorNmos: 1.89207e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.42146e+08 muA
** DiodeTransistorPmos: -6.37209e+07 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** inputVoltageBiasXXpXX2: 4.26201  V
** out: 2.5  V
** outFirstStage: 4.03701  V
** outVoltageBiasXXnXX1: 1.09701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.700001  V
** innerStageBias: 0.542001  V
** out1: 1.32301  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.60101  V


.END